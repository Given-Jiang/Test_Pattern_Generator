-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.1.0 Build 162 10/23/2013 SJ Full Version
-- Created on Wed Feb 11 10:18:10 2015

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY StateMachineEditor1 IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        col_select : IN STD_LOGIC_VECTOR(2 DOWNTO 0) := "000";
        data_en : IN STD_LOGIC := '0';
        data : OUT STD_LOGIC_VECTOR(23 DOWNTO 0)
    );
END StateMachineEditor1;

ARCHITECTURE BEHAVIOR OF StateMachineEditor1 IS
    TYPE type_fstate IS (IDLE,BLOCKA,BLOCKB,BLOCKC);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,col_select,data_en)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= IDLE;
            data <= "000000000000000000000000";
        ELSE
            data <= "000000000000000000000000";
            CASE fstate IS
                WHEN IDLE =>
                    IF (((col_select(2 DOWNTO 0) = "001") AND (data_en = '1'))) THEN
                        reg_fstate <= BLOCKA;
                    ELSIF ((col_select(2 DOWNTO 0) = "000")) THEN
                        reg_fstate <= IDLE;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= IDLE;
                    END IF;

                    data <= "000000000000000000000000";
                WHEN BLOCKA =>
                    IF (((col_select(2 DOWNTO 0) = "010") AND (data_en = '1'))) THEN
                        reg_fstate <= BLOCKB;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= BLOCKA;
                    END IF;

                    data <= "000000000000000011111111";
                WHEN BLOCKB =>
                    IF (((col_select(2 DOWNTO 0) = "100") AND (data_en = '1'))) THEN
                        reg_fstate <= BLOCKC;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= BLOCKB;
                    END IF;

                    data <= "000000001111111100000000";
                WHEN BLOCKC =>
                    IF ((col_select(2 DOWNTO 0) = "000")) THEN
                        reg_fstate <= IDLE;
                    ELSIF (((col_select(2 DOWNTO 0) = "001") AND (data_en = '1'))) THEN
                        reg_fstate <= BLOCKA;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= BLOCKC;
                    END IF;

                    data <= "111111110000000000000000";
                WHEN OTHERS => 
                    data <= "XXXXXXXXXXXXXXXXXXXXXXXX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
