-- Test_Pattern_Generator_GN_Test_Pattern_Generator_CTRL_PAK_TRANSLATE.vhd

-- Generated using ACDS version 13.1 162 at 2015.02.27.10:05:29

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Test_Pattern_Generator_GN_Test_Pattern_Generator_CTRL_PAK_TRANSLATE is
	port (
		ctrl_pak2 : out std_logic_vector(23 downto 0);                    -- ctrl_pak2.wire
		dil       : in  std_logic_vector(3 downto 0)  := (others => '0'); --       dil.wire
		col       : in  std_logic_vector(31 downto 0) := (others => '0'); --       col.wire
		Clock     : in  std_logic                     := '0';             --     Clock.clk
		aclr      : in  std_logic                     := '0';             --          .reset
		ctrl_pak1 : out std_logic_vector(23 downto 0);                    -- ctrl_pak1.wire
		ctrl_pak3 : out std_logic_vector(23 downto 0);                    -- ctrl_pak3.wire
		row       : in  std_logic_vector(31 downto 0) := (others => '0')  --       row.wire
	);
end entity Test_Pattern_Generator_GN_Test_Pattern_Generator_CTRL_PAK_TRANSLATE;

architecture rtl of Test_Pattern_Generator_GN_Test_Pattern_Generator_CTRL_PAK_TRANSLATE is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_cast_GNTS3MQUMJ is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(3 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GNTS3MQUMJ;

	component alt_dspbuilder_port_GNEPKLLZKY is
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNEPKLLZKY;

	component alt_dspbuilder_cast_GNJ7VFHJ4A is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(3 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GNJ7VFHJ4A;

	component alt_dspbuilder_cast_GNMYKU6OLE is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(3 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GNMYKU6OLE;

	component alt_dspbuilder_cast_GN5VN2FCXZ is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(3 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GN5VN2FCXZ;

	component alt_dspbuilder_bus_concat_GNAUBM7IRL is
		generic (
			widthB : natural := 8;
			widthA : natural := 8
		);
		port (
			a      : in  std_logic_vector(widthA-1 downto 0)        := (others => 'X'); -- wire
			aclr   : in  std_logic                                  := 'X';             -- clk
			b      : in  std_logic_vector(widthB-1 downto 0)        := (others => 'X'); -- wire
			clock  : in  std_logic                                  := 'X';             -- clk
			output : out std_logic_vector(widthA+widthB-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_bus_concat_GNAUBM7IRL;

	component alt_dspbuilder_bus_concat_GNWZPLIVXS is
		generic (
			widthB : natural := 8;
			widthA : natural := 8
		);
		port (
			a      : in  std_logic_vector(widthA-1 downto 0)        := (others => 'X'); -- wire
			aclr   : in  std_logic                                  := 'X';             -- clk
			b      : in  std_logic_vector(widthB-1 downto 0)        := (others => 'X'); -- wire
			clock  : in  std_logic                                  := 'X';             -- clk
			output : out std_logic_vector(widthA+widthB-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_bus_concat_GNWZPLIVXS;

	component alt_dspbuilder_bus_concat_GNIIOZRPJD is
		generic (
			widthB : natural := 8;
			widthA : natural := 8
		);
		port (
			a      : in  std_logic_vector(widthA-1 downto 0)        := (others => 'X'); -- wire
			aclr   : in  std_logic                                  := 'X';             -- clk
			b      : in  std_logic_vector(widthB-1 downto 0)        := (others => 'X'); -- wire
			clock  : in  std_logic                                  := 'X';             -- clk
			output : out std_logic_vector(widthA+widthB-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_bus_concat_GNIIOZRPJD;

	component alt_dspbuilder_port_GNOC3SGKQJ is
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNOC3SGKQJ;

	component alt_dspbuilder_constant_GNPLBTTHPL is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(3 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNPLBTTHPL;

	component alt_dspbuilder_port_GNCNBVQF75 is
		port (
			input  : in  std_logic_vector(3 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(3 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNCNBVQF75;

	component alt_dspbuilder_bus_concat_GN55ETJ4VI is
		generic (
			widthB : natural := 8;
			widthA : natural := 8
		);
		port (
			a      : in  std_logic_vector(widthA-1 downto 0)        := (others => 'X'); -- wire
			aclr   : in  std_logic                                  := 'X';             -- clk
			b      : in  std_logic_vector(widthB-1 downto 0)        := (others => 'X'); -- wire
			clock  : in  std_logic                                  := 'X';             -- clk
			output : out std_logic_vector(widthA+widthB-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_bus_concat_GN55ETJ4VI;

	component alt_dspbuilder_cast_GNMMXHT3UH is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(3 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(3 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNMMXHT3UH;

	component alt_dspbuilder_cast_GNNZHXLS76 is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(15 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNNZHXLS76;

	signal bus_concatenation12_output_wire : std_logic_vector(15 downto 0); -- Bus_Concatenation12:output -> Bus_Concatenation13:a
	signal bus_concatenation10_output_wire : std_logic_vector(7 downto 0);  -- Bus_Concatenation10:output -> Bus_Concatenation14:a
	signal bus_concatenation11_output_wire : std_logic_vector(7 downto 0);  -- Bus_Concatenation11:output -> Bus_Concatenation14:b
	signal bus_concatenation15_output_wire : std_logic_vector(7 downto 0);  -- Bus_Concatenation15:output -> Bus_Concatenation16:a
	signal bus_concatenation14_output_wire : std_logic_vector(15 downto 0); -- Bus_Concatenation14:output -> Bus_Concatenation16:b
	signal bus_concatenation5_output_wire  : std_logic_vector(7 downto 0);  -- Bus_Concatenation5:output -> Bus_Concatenation13:b
	signal bus_concatenation2_output_wire  : std_logic_vector(7 downto 0);  -- Bus_Concatenation2:output -> Bus_Concatenation6:a
	signal bus_concatenation3_output_wire  : std_logic_vector(7 downto 0);  -- Bus_Concatenation3:output -> Bus_Concatenation6:b
	signal bus_concatenation7_output_wire  : std_logic_vector(7 downto 0);  -- Bus_Concatenation7:output -> Bus_Concatenation12:a
	signal bus_concatenation6_output_wire  : std_logic_vector(15 downto 0); -- Bus_Concatenation6:output -> Bus_Concatenation8:a
	signal bus_concatenation4_output_wire  : std_logic_vector(7 downto 0);  -- Bus_Concatenation4:output -> Bus_Concatenation8:b
	signal bus_concatenation9_output_wire  : std_logic_vector(7 downto 0);  -- Bus_Concatenation9:output -> Bus_Concatenation12:b
	signal bus_conversion_output_wire      : std_logic_vector(3 downto 0);  -- Bus_Conversion:output -> Bus_Concatenation3:b
	signal bus_conversion2_output_wire     : std_logic_vector(3 downto 0);  -- Bus_Conversion2:output -> Bus_Concatenation2:b
	signal bus_conversion3_output_wire     : std_logic_vector(3 downto 0);  -- Bus_Conversion3:output -> Bus_Concatenation5:b
	signal bus_conversion4_output_wire     : std_logic_vector(3 downto 0);  -- Bus_Conversion4:output -> Bus_Concatenation4:b
	signal bus_conversion5_output_wire     : std_logic_vector(3 downto 0);  -- Bus_Conversion5:output -> Bus_Concatenation9:b
	signal bus_conversion6_output_wire     : std_logic_vector(3 downto 0);  -- Bus_Conversion6:output -> Bus_Concatenation7:b
	signal bus_conversion7_output_wire     : std_logic_vector(3 downto 0);  -- Bus_Conversion7:output -> Bus_Concatenation11:b
	signal bus_conversion8_output_wire     : std_logic_vector(3 downto 0);  -- Bus_Conversion8:output -> Bus_Concatenation10:b
	signal bus_concatenation8_output_wire  : std_logic_vector(23 downto 0); -- Bus_Concatenation8:output -> ctrl_pak1_0:input
	signal bus_concatenation13_output_wire : std_logic_vector(23 downto 0); -- Bus_Concatenation13:output -> ctrl_pak2_0:input
	signal bus_concatenation16_output_wire : std_logic_vector(23 downto 0); -- Bus_Concatenation16:output -> ctrl_pak3_0:input
	signal dil_0_output_wire               : std_logic_vector(3 downto 0);  -- dil_0:output -> cast8:input
	signal cast8_output_wire               : std_logic_vector(3 downto 0);  -- cast8:output -> Bus_Concatenation15:b
	signal col_0_output_wire               : std_logic_vector(31 downto 0); -- col_0:output -> [cast10:input, cast11:input, cast12:input, cast9:input]
	signal cast9_output_wire               : std_logic_vector(15 downto 0); -- cast9:output -> Bus_Conversion:input
	signal cast10_output_wire              : std_logic_vector(15 downto 0); -- cast10:output -> Bus_Conversion2:input
	signal cast11_output_wire              : std_logic_vector(15 downto 0); -- cast11:output -> Bus_Conversion3:input
	signal cast12_output_wire              : std_logic_vector(15 downto 0); -- cast12:output -> Bus_Conversion4:input
	signal row_0_output_wire               : std_logic_vector(31 downto 0); -- row_0:output -> [cast13:input, cast14:input, cast15:input, cast16:input]
	signal cast13_output_wire              : std_logic_vector(15 downto 0); -- cast13:output -> Bus_Conversion5:input
	signal cast14_output_wire              : std_logic_vector(15 downto 0); -- cast14:output -> Bus_Conversion6:input
	signal cast15_output_wire              : std_logic_vector(15 downto 0); -- cast15:output -> Bus_Conversion7:input
	signal cast16_output_wire              : std_logic_vector(15 downto 0); -- cast16:output -> Bus_Conversion8:input
	signal constant10_output_wire          : std_logic_vector(3 downto 0);  -- Constant10:output -> cast17:input
	signal cast17_output_wire              : std_logic_vector(3 downto 0);  -- cast17:output -> Bus_Concatenation2:a
	signal constant19_output_wire          : std_logic_vector(3 downto 0);  -- Constant19:output -> cast18:input
	signal cast18_output_wire              : std_logic_vector(3 downto 0);  -- cast18:output -> Bus_Concatenation3:a
	signal constant21_output_wire          : std_logic_vector(3 downto 0);  -- Constant21:output -> cast19:input
	signal cast19_output_wire              : std_logic_vector(3 downto 0);  -- cast19:output -> Bus_Concatenation4:a
	signal constant22_output_wire          : std_logic_vector(3 downto 0);  -- Constant22:output -> cast20:input
	signal cast20_output_wire              : std_logic_vector(3 downto 0);  -- cast20:output -> Bus_Concatenation5:a
	signal constant23_output_wire          : std_logic_vector(3 downto 0);  -- Constant23:output -> cast21:input
	signal cast21_output_wire              : std_logic_vector(3 downto 0);  -- cast21:output -> Bus_Concatenation7:a
	signal constant24_output_wire          : std_logic_vector(3 downto 0);  -- Constant24:output -> cast22:input
	signal cast22_output_wire              : std_logic_vector(3 downto 0);  -- cast22:output -> Bus_Concatenation9:a
	signal constant25_output_wire          : std_logic_vector(3 downto 0);  -- Constant25:output -> cast23:input
	signal cast23_output_wire              : std_logic_vector(3 downto 0);  -- cast23:output -> Bus_Concatenation10:a
	signal constant26_output_wire          : std_logic_vector(3 downto 0);  -- Constant26:output -> cast24:input
	signal cast24_output_wire              : std_logic_vector(3 downto 0);  -- cast24:output -> Bus_Concatenation11:a
	signal constant27_output_wire          : std_logic_vector(3 downto 0);  -- Constant27:output -> cast25:input
	signal cast25_output_wire              : std_logic_vector(3 downto 0);  -- cast25:output -> Bus_Concatenation15:a
	signal clock_0_clock_output_reset      : std_logic;                     -- Clock_0:aclr_out -> [Bus_Concatenation10:aclr, Bus_Concatenation11:aclr, Bus_Concatenation12:aclr, Bus_Concatenation13:aclr, Bus_Concatenation14:aclr, Bus_Concatenation15:aclr, Bus_Concatenation16:aclr, Bus_Concatenation2:aclr, Bus_Concatenation3:aclr, Bus_Concatenation4:aclr, Bus_Concatenation5:aclr, Bus_Concatenation6:aclr, Bus_Concatenation7:aclr, Bus_Concatenation8:aclr, Bus_Concatenation9:aclr]
	signal clock_0_clock_output_clk        : std_logic;                     -- Clock_0:clock_out -> [Bus_Concatenation10:clock, Bus_Concatenation11:clock, Bus_Concatenation12:clock, Bus_Concatenation13:clock, Bus_Concatenation14:clock, Bus_Concatenation15:clock, Bus_Concatenation16:clock, Bus_Concatenation2:clock, Bus_Concatenation3:clock, Bus_Concatenation4:clock, Bus_Concatenation5:clock, Bus_Concatenation6:clock, Bus_Concatenation7:clock, Bus_Concatenation8:clock, Bus_Concatenation9:clock]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	bus_conversion2 : component alt_dspbuilder_cast_GNTS3MQUMJ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast10_output_wire,          --  input.wire
			output => bus_conversion2_output_wire  -- output.wire
		);

	col_0 : component alt_dspbuilder_port_GNEPKLLZKY
		port map (
			input  => col,               --  input.wire
			output => col_0_output_wire  -- output.wire
		);

	bus_conversion3 : component alt_dspbuilder_cast_GNJ7VFHJ4A
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast11_output_wire,          --  input.wire
			output => bus_conversion3_output_wire  -- output.wire
		);

	bus_conversion4 : component alt_dspbuilder_cast_GNMYKU6OLE
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast12_output_wire,          --  input.wire
			output => bus_conversion4_output_wire  -- output.wire
		);

	bus_conversion : component alt_dspbuilder_cast_GN5VN2FCXZ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast9_output_wire,          --  input.wire
			output => bus_conversion_output_wire  -- output.wire
		);

	bus_concatenation7 : component alt_dspbuilder_bus_concat_GNAUBM7IRL
		generic map (
			widthB => 4,
			widthA => 4
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => cast21_output_wire,             --          a.wire
			b      => bus_conversion6_output_wire,    --          b.wire
			output => bus_concatenation7_output_wire  --     output.wire
		);

	bus_concatenation8 : component alt_dspbuilder_bus_concat_GNWZPLIVXS
		generic map (
			widthB => 8,
			widthA => 16
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => bus_concatenation6_output_wire, --          a.wire
			b      => bus_concatenation4_output_wire, --          b.wire
			output => bus_concatenation8_output_wire  --     output.wire
		);

	bus_concatenation5 : component alt_dspbuilder_bus_concat_GNAUBM7IRL
		generic map (
			widthB => 4,
			widthA => 4
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => cast20_output_wire,             --          a.wire
			b      => bus_conversion3_output_wire,    --          b.wire
			output => bus_concatenation5_output_wire  --     output.wire
		);

	bus_concatenation6 : component alt_dspbuilder_bus_concat_GNIIOZRPJD
		generic map (
			widthB => 8,
			widthA => 8
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => bus_concatenation2_output_wire, --          a.wire
			b      => bus_concatenation3_output_wire, --          b.wire
			output => bus_concatenation6_output_wire  --     output.wire
		);

	bus_concatenation3 : component alt_dspbuilder_bus_concat_GNAUBM7IRL
		generic map (
			widthB => 4,
			widthA => 4
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => cast18_output_wire,             --          a.wire
			b      => bus_conversion_output_wire,     --          b.wire
			output => bus_concatenation3_output_wire  --     output.wire
		);

	bus_concatenation4 : component alt_dspbuilder_bus_concat_GNAUBM7IRL
		generic map (
			widthB => 4,
			widthA => 4
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => cast19_output_wire,             --          a.wire
			b      => bus_conversion4_output_wire,    --          b.wire
			output => bus_concatenation4_output_wire  --     output.wire
		);

	bus_concatenation2 : component alt_dspbuilder_bus_concat_GNAUBM7IRL
		generic map (
			widthB => 4,
			widthA => 4
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => cast17_output_wire,             --          a.wire
			b      => bus_conversion2_output_wire,    --          b.wire
			output => bus_concatenation2_output_wire  --     output.wire
		);

	ctrl_pak2_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => bus_concatenation13_output_wire, --  input.wire
			output => ctrl_pak2                        -- output.wire
		);

	ctrl_pak3_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => bus_concatenation16_output_wire, --  input.wire
			output => ctrl_pak3                        -- output.wire
		);

	constant10 : component alt_dspbuilder_constant_GNPLBTTHPL
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "0000",
			width      => 4
		)
		port map (
			output => constant10_output_wire  -- output.wire
		);

	ctrl_pak1_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => bus_concatenation8_output_wire, --  input.wire
			output => ctrl_pak1                       -- output.wire
		);

	constant19 : component alt_dspbuilder_constant_GNPLBTTHPL
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "0000",
			width      => 4
		)
		port map (
			output => constant19_output_wire  -- output.wire
		);

	dil_0 : component alt_dspbuilder_port_GNCNBVQF75
		port map (
			input  => dil,               --  input.wire
			output => dil_0_output_wire  -- output.wire
		);

	constant27 : component alt_dspbuilder_constant_GNPLBTTHPL
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "0000",
			width      => 4
		)
		port map (
			output => constant27_output_wire  -- output.wire
		);

	constant26 : component alt_dspbuilder_constant_GNPLBTTHPL
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "0000",
			width      => 4
		)
		port map (
			output => constant26_output_wire  -- output.wire
		);

	constant23 : component alt_dspbuilder_constant_GNPLBTTHPL
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "0000",
			width      => 4
		)
		port map (
			output => constant23_output_wire  -- output.wire
		);

	bus_concatenation13 : component alt_dspbuilder_bus_concat_GNWZPLIVXS
		generic map (
			widthB => 8,
			widthA => 16
		)
		port map (
			clock  => clock_0_clock_output_clk,        -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,      --           .reset
			a      => bus_concatenation12_output_wire, --          a.wire
			b      => bus_concatenation5_output_wire,  --          b.wire
			output => bus_concatenation13_output_wire  --     output.wire
		);

	constant22 : component alt_dspbuilder_constant_GNPLBTTHPL
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "0000",
			width      => 4
		)
		port map (
			output => constant22_output_wire  -- output.wire
		);

	bus_concatenation12 : component alt_dspbuilder_bus_concat_GNIIOZRPJD
		generic map (
			widthB => 8,
			widthA => 8
		)
		port map (
			clock  => clock_0_clock_output_clk,        -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,      --           .reset
			a      => bus_concatenation7_output_wire,  --          a.wire
			b      => bus_concatenation9_output_wire,  --          b.wire
			output => bus_concatenation12_output_wire  --     output.wire
		);

	constant25 : component alt_dspbuilder_constant_GNPLBTTHPL
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "0000",
			width      => 4
		)
		port map (
			output => constant25_output_wire  -- output.wire
		);

	bus_concatenation11 : component alt_dspbuilder_bus_concat_GNAUBM7IRL
		generic map (
			widthB => 4,
			widthA => 4
		)
		port map (
			clock  => clock_0_clock_output_clk,        -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,      --           .reset
			a      => cast24_output_wire,              --          a.wire
			b      => bus_conversion7_output_wire,     --          b.wire
			output => bus_concatenation11_output_wire  --     output.wire
		);

	constant24 : component alt_dspbuilder_constant_GNPLBTTHPL
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "0000",
			width      => 4
		)
		port map (
			output => constant24_output_wire  -- output.wire
		);

	bus_concatenation10 : component alt_dspbuilder_bus_concat_GNAUBM7IRL
		generic map (
			widthB => 4,
			widthA => 4
		)
		port map (
			clock  => clock_0_clock_output_clk,        -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,      --           .reset
			a      => cast23_output_wire,              --          a.wire
			b      => bus_conversion8_output_wire,     --          b.wire
			output => bus_concatenation10_output_wire  --     output.wire
		);

	bus_concatenation16 : component alt_dspbuilder_bus_concat_GN55ETJ4VI
		generic map (
			widthB => 16,
			widthA => 8
		)
		port map (
			clock  => clock_0_clock_output_clk,        -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,      --           .reset
			a      => bus_concatenation15_output_wire, --          a.wire
			b      => bus_concatenation14_output_wire, --          b.wire
			output => bus_concatenation16_output_wire  --     output.wire
		);

	constant21 : component alt_dspbuilder_constant_GNPLBTTHPL
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "0000",
			width      => 4
		)
		port map (
			output => constant21_output_wire  -- output.wire
		);

	bus_concatenation15 : component alt_dspbuilder_bus_concat_GNAUBM7IRL
		generic map (
			widthB => 4,
			widthA => 4
		)
		port map (
			clock  => clock_0_clock_output_clk,        -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,      --           .reset
			a      => cast25_output_wire,              --          a.wire
			b      => cast8_output_wire,               --          b.wire
			output => bus_concatenation15_output_wire  --     output.wire
		);

	row_0 : component alt_dspbuilder_port_GNEPKLLZKY
		port map (
			input  => row,               --  input.wire
			output => row_0_output_wire  -- output.wire
		);

	bus_concatenation14 : component alt_dspbuilder_bus_concat_GNIIOZRPJD
		generic map (
			widthB => 8,
			widthA => 8
		)
		port map (
			clock  => clock_0_clock_output_clk,        -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,      --           .reset
			a      => bus_concatenation10_output_wire, --          a.wire
			b      => bus_concatenation11_output_wire, --          b.wire
			output => bus_concatenation14_output_wire  --     output.wire
		);

	bus_concatenation9 : component alt_dspbuilder_bus_concat_GNAUBM7IRL
		generic map (
			widthB => 4,
			widthA => 4
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => cast22_output_wire,             --          a.wire
			b      => bus_conversion5_output_wire,    --          b.wire
			output => bus_concatenation9_output_wire  --     output.wire
		);

	bus_conversion8 : component alt_dspbuilder_cast_GNJ7VFHJ4A
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast16_output_wire,          --  input.wire
			output => bus_conversion8_output_wire  -- output.wire
		);

	bus_conversion7 : component alt_dspbuilder_cast_GNTS3MQUMJ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast15_output_wire,          --  input.wire
			output => bus_conversion7_output_wire  -- output.wire
		);

	bus_conversion6 : component alt_dspbuilder_cast_GN5VN2FCXZ
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast14_output_wire,          --  input.wire
			output => bus_conversion6_output_wire  -- output.wire
		);

	bus_conversion5 : component alt_dspbuilder_cast_GNMYKU6OLE
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => cast13_output_wire,          --  input.wire
			output => bus_conversion5_output_wire  -- output.wire
		);

	cast8 : component alt_dspbuilder_cast_GNMMXHT3UH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => dil_0_output_wire, --  input.wire
			output => cast8_output_wire  -- output.wire
		);

	cast9 : component alt_dspbuilder_cast_GNNZHXLS76
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => col_0_output_wire, --  input.wire
			output => cast9_output_wire  -- output.wire
		);

	cast10 : component alt_dspbuilder_cast_GNNZHXLS76
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => col_0_output_wire,  --  input.wire
			output => cast10_output_wire  -- output.wire
		);

	cast11 : component alt_dspbuilder_cast_GNNZHXLS76
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => col_0_output_wire,  --  input.wire
			output => cast11_output_wire  -- output.wire
		);

	cast12 : component alt_dspbuilder_cast_GNNZHXLS76
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => col_0_output_wire,  --  input.wire
			output => cast12_output_wire  -- output.wire
		);

	cast13 : component alt_dspbuilder_cast_GNNZHXLS76
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => row_0_output_wire,  --  input.wire
			output => cast13_output_wire  -- output.wire
		);

	cast14 : component alt_dspbuilder_cast_GNNZHXLS76
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => row_0_output_wire,  --  input.wire
			output => cast14_output_wire  -- output.wire
		);

	cast15 : component alt_dspbuilder_cast_GNNZHXLS76
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => row_0_output_wire,  --  input.wire
			output => cast15_output_wire  -- output.wire
		);

	cast16 : component alt_dspbuilder_cast_GNNZHXLS76
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => row_0_output_wire,  --  input.wire
			output => cast16_output_wire  -- output.wire
		);

	cast17 : component alt_dspbuilder_cast_GNMMXHT3UH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant10_output_wire, --  input.wire
			output => cast17_output_wire      -- output.wire
		);

	cast18 : component alt_dspbuilder_cast_GNMMXHT3UH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant19_output_wire, --  input.wire
			output => cast18_output_wire      -- output.wire
		);

	cast19 : component alt_dspbuilder_cast_GNMMXHT3UH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant21_output_wire, --  input.wire
			output => cast19_output_wire      -- output.wire
		);

	cast20 : component alt_dspbuilder_cast_GNMMXHT3UH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant22_output_wire, --  input.wire
			output => cast20_output_wire      -- output.wire
		);

	cast21 : component alt_dspbuilder_cast_GNMMXHT3UH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant23_output_wire, --  input.wire
			output => cast21_output_wire      -- output.wire
		);

	cast22 : component alt_dspbuilder_cast_GNMMXHT3UH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant24_output_wire, --  input.wire
			output => cast22_output_wire      -- output.wire
		);

	cast23 : component alt_dspbuilder_cast_GNMMXHT3UH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant25_output_wire, --  input.wire
			output => cast23_output_wire      -- output.wire
		);

	cast24 : component alt_dspbuilder_cast_GNMMXHT3UH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant26_output_wire, --  input.wire
			output => cast24_output_wire      -- output.wire
		);

	cast25 : component alt_dspbuilder_cast_GNMMXHT3UH
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant27_output_wire, --  input.wire
			output => cast25_output_wire      -- output.wire
		);

end architecture rtl; -- of Test_Pattern_Generator_GN_Test_Pattern_Generator_CTRL_PAK_TRANSLATE
