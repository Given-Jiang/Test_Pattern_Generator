-- Test_Pattern_Generator_GN.vhd

-- Generated using ACDS version 13.1 162 at 2015.02.27.10:05:29

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Test_Pattern_Generator_GN is
	port (
		Clock                          : in  std_logic                     := '0';             --                          Clock.clk
		aclr                           : in  std_logic                     := '0';             --                               .reset_n
		Avalon_ST_Source_ready         : in  std_logic                     := '0';             --         Avalon_ST_Source_ready.wire
		Avalon_ST_Source_valid         : out std_logic;                                        --         Avalon_ST_Source_valid.wire
		Avalon_MM_Slave_write          : in  std_logic                     := '0';             --          Avalon_MM_Slave_write.wire
		Avalon_MM_Slave_writedata      : in  std_logic_vector(31 downto 0) := (others => '0'); --      Avalon_MM_Slave_writedata.wire
		Avalon_ST_Source_endofpacket   : out std_logic;                                        --   Avalon_ST_Source_endofpacket.wire
		Avalon_ST_Source_data          : out std_logic_vector(23 downto 0);                    --          Avalon_ST_Source_data.wire
		Avalon_MM_Slave_address        : in  std_logic_vector(1 downto 0)  := (others => '0'); --        Avalon_MM_Slave_address.wire
		Avalon_ST_Source_startofpacket : out std_logic                                         -- Avalon_ST_Source_startofpacket.wire
	);
end entity Test_Pattern_Generator_GN;

architecture rtl of Test_Pattern_Generator_GN is
	component alt_dspbuilder_clock_GNF343OQUJ is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNF343OQUJ;

	component alt_dspbuilder_port_GN6TDLHAW6 is
		port (
			input  : in  std_logic_vector(1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GN6TDLHAW6;

	component Test_Pattern_Generator_GN_Test_Pattern_Generator_DATA_GENERATE is
		port (
			Clock    : in  std_logic                     := 'X';             -- clk
			aclr     : in  std_logic                     := 'X';             -- reset
			counter  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			col      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			colorbar : out std_logic_vector(23 downto 0);                    -- wire
			data_en  : in  std_logic                     := 'X';             -- wire
			ctrl_en  : in  std_logic                     := 'X'              -- wire
		);
	end component Test_Pattern_Generator_GN_Test_Pattern_Generator_DATA_GENERATE;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_port_GNEPKLLZKY is
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNEPKLLZKY;

	component Test_Pattern_Generator_GN_Test_Pattern_Generator_CTRL_PAK_TRANSLATE is
		port (
			ctrl_pak2 : out std_logic_vector(23 downto 0);                    -- wire
			dil       : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- wire
			col       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			Clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			ctrl_pak1 : out std_logic_vector(23 downto 0);                    -- wire
			ctrl_pak3 : out std_logic_vector(23 downto 0);                    -- wire
			row       : in  std_logic_vector(31 downto 0) := (others => 'X')  -- wire
		);
	end component Test_Pattern_Generator_GN_Test_Pattern_Generator_CTRL_PAK_TRANSLATE;

	component alt_dspbuilder_constant_GNPLBTTHPL is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(3 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNPLBTTHPL;

	component alt_dspbuilder_delay_GNPJ4Y7BVC is
		generic (
			ClockPhase : string   := "1";
			delay      : positive := 1;
			use_init   : natural  := 0;
			BitPattern : string   := "00000001";
			width      : positive := 8
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNPJ4Y7BVC;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_logical_bit_op_GNUQ2R64DV is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'; -- wire
			data1  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNUQ2R64DV;

	component alt_dspbuilder_port_GNOC3SGKQJ is
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNOC3SGKQJ;

	component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'; -- wire
			data1  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V;

	component alt_dspbuilder_decoder_GNEQGKKPXW is
		generic (
			decode   : string  := "00000000";
			pipeline : natural := 0;
			width    : natural := 8
		);
		port (
			aclr  : in  std_logic                          := 'X';             -- clk
			clock : in  std_logic                          := 'X';             -- clk
			data  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			dec   : out std_logic;                                             -- wire
			ena   : in  std_logic                          := 'X';             -- wire
			sclr  : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_decoder_GNEQGKKPXW;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component Test_Pattern_Generator_GN_Test_Pattern_Generator_MAIN_CTRL is
		port (
			eop       : out std_logic;                                        -- wire
			counter_1 : out std_logic_vector(23 downto 0);                    -- wire
			colorbar  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			data      : out std_logic_vector(24 downto 0);                    -- wire
			col       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			ctrl_pak3 : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			ctrl_pak2 : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			data_en   : out std_logic;                                        -- wire
			ctrl_en   : out std_logic;                                        -- wire
			Clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			row       : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			ctrl_pak1 : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			check_en  : out std_logic;                                        -- wire
			sop       : out std_logic;                                        -- wire
			ready     : in  std_logic                     := 'X'              -- wire
		);
	end component Test_Pattern_Generator_GN_Test_Pattern_Generator_MAIN_CTRL;

	component alt_dspbuilder_decoder_GNM4LOIHXZ is
		generic (
			decode   : string  := "00000000";
			pipeline : natural := 0;
			width    : natural := 8
		);
		port (
			aclr  : in  std_logic                          := 'X';             -- clk
			clock : in  std_logic                          := 'X';             -- clk
			data  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			dec   : out std_logic;                                             -- wire
			ena   : in  std_logic                          := 'X';             -- wire
			sclr  : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_decoder_GNM4LOIHXZ;

	component alt_dspbuilder_cast_GN5EYRLJQW is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(24 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN5EYRLJQW;

	signal delaysclrgnd_output_wire                                   : std_logic;                     -- DelaysclrGND:output -> Delay:sclr
	signal decoder1sclrgnd_output_wire                                : std_logic;                     -- Decoder1sclrGND:output -> Decoder1:sclr
	signal decoder1enavcc_output_wire                                 : std_logic;                     -- Decoder1enaVCC:output -> Decoder1:ena
	signal delay3sclrgnd_output_wire                                  : std_logic;                     -- Delay3sclrGND:output -> Delay3:sclr
	signal delay1sclrgnd_output_wire                                  : std_logic;                     -- Delay1sclrGND:output -> Delay1:sclr
	signal delay2sclrgnd_output_wire                                  : std_logic;                     -- Delay2sclrGND:output -> Delay2:sclr
	signal decodersclrgnd_output_wire                                 : std_logic;                     -- DecodersclrGND:output -> Decoder:sclr
	signal decoderenavcc_output_wire                                  : std_logic;                     -- DecoderenaVCC:output -> Decoder:ena
	signal avalon_mm_slave_address_0_output_wire                      : std_logic_vector(1 downto 0);  -- Avalon_MM_Slave_address_0:output -> [Decoder1:data, Decoder:data]
	signal delay_output_wire                                          : std_logic_vector(31 downto 0); -- Delay:output -> Delay2:input
	signal delay1_output_wire                                         : std_logic_vector(31 downto 0); -- Delay1:output -> Delay3:input
	signal constant3_output_wire                                      : std_logic_vector(3 downto 0);  -- Constant3:output -> Test_Pattern_Generator_CTRL_PAK_TRANSLATE_0:dil
	signal delay2_output_wire                                         : std_logic_vector(31 downto 0); -- Delay2:output -> [Test_Pattern_Generator_CTRL_PAK_TRANSLATE_0:col, Test_Pattern_Generator_DATA_GENERATE_0:col, Test_Pattern_Generator_MAIN_CTRL_0:col]
	signal delay3_output_wire                                         : std_logic_vector(31 downto 0); -- Delay3:output -> [Test_Pattern_Generator_CTRL_PAK_TRANSLATE_0:row, Test_Pattern_Generator_MAIN_CTRL_0:row]
	signal avalon_mm_slave_writedata_0_output_wire                    : std_logic_vector(31 downto 0); -- Avalon_MM_Slave_writedata_0:output -> [Delay1:input, Delay:input]
	signal test_pattern_generator_main_ctrl_0_check_en_wire           : std_logic;                     -- Test_Pattern_Generator_MAIN_CTRL_0:check_en -> [Delay2:ena, Delay3:ena]
	signal decoder_dec_wire                                           : std_logic;                     -- Decoder:dec -> Logical_Bit_Operator:data0
	signal avalon_mm_slave_write_0_output_wire                        : std_logic;                     -- Avalon_MM_Slave_write_0:output -> [Logical_Bit_Operator1:data0, Logical_Bit_Operator:data1]
	signal logical_bit_operator_result_wire                           : std_logic;                     -- Logical_Bit_Operator:result -> Delay:ena
	signal decoder1_dec_wire                                          : std_logic;                     -- Decoder1:dec -> Logical_Bit_Operator1:data1
	signal logical_bit_operator1_result_wire                          : std_logic;                     -- Logical_Bit_Operator1:result -> Delay1:ena
	signal logical_bit_operator2_result_wire                          : std_logic;                     -- Logical_Bit_Operator2:result -> Avalon_ST_Source_valid_0:input
	signal avalon_st_source_ready_0_output_wire                       : std_logic;                     -- Avalon_ST_Source_ready_0:output -> Test_Pattern_Generator_MAIN_CTRL_0:ready
	signal test_pattern_generator_ctrl_pak_translate_0_ctrl_pak1_wire : std_logic_vector(23 downto 0); -- Test_Pattern_Generator_CTRL_PAK_TRANSLATE_0:ctrl_pak1 -> Test_Pattern_Generator_MAIN_CTRL_0:ctrl_pak1
	signal test_pattern_generator_ctrl_pak_translate_0_ctrl_pak2_wire : std_logic_vector(23 downto 0); -- Test_Pattern_Generator_CTRL_PAK_TRANSLATE_0:ctrl_pak2 -> Test_Pattern_Generator_MAIN_CTRL_0:ctrl_pak2
	signal test_pattern_generator_ctrl_pak_translate_0_ctrl_pak3_wire : std_logic_vector(23 downto 0); -- Test_Pattern_Generator_CTRL_PAK_TRANSLATE_0:ctrl_pak3 -> Test_Pattern_Generator_MAIN_CTRL_0:ctrl_pak3
	signal test_pattern_generator_data_generate_0_colorbar_wire       : std_logic_vector(23 downto 0); -- Test_Pattern_Generator_DATA_GENERATE_0:colorbar -> Test_Pattern_Generator_MAIN_CTRL_0:colorbar
	signal test_pattern_generator_main_ctrl_0_ctrl_en_wire            : std_logic;                     -- Test_Pattern_Generator_MAIN_CTRL_0:ctrl_en -> [Logical_Bit_Operator2:data0, Test_Pattern_Generator_DATA_GENERATE_0:ctrl_en]
	signal test_pattern_generator_main_ctrl_0_data_en_wire            : std_logic;                     -- Test_Pattern_Generator_MAIN_CTRL_0:data_en -> [Logical_Bit_Operator2:data1, Test_Pattern_Generator_DATA_GENERATE_0:data_en]
	signal test_pattern_generator_main_ctrl_0_sop_wire                : std_logic;                     -- Test_Pattern_Generator_MAIN_CTRL_0:sop -> Avalon_ST_Source_startofpacket_0:input
	signal test_pattern_generator_main_ctrl_0_eop_wire                : std_logic;                     -- Test_Pattern_Generator_MAIN_CTRL_0:eop -> Avalon_ST_Source_endofpacket_0:input
	signal test_pattern_generator_main_ctrl_0_counter_1_wire          : std_logic_vector(23 downto 0); -- Test_Pattern_Generator_MAIN_CTRL_0:counter_1 -> Test_Pattern_Generator_DATA_GENERATE_0:counter
	signal test_pattern_generator_main_ctrl_0_data_wire               : std_logic_vector(24 downto 0); -- Test_Pattern_Generator_MAIN_CTRL_0:data -> cast44:input
	signal cast44_output_wire                                         : std_logic_vector(23 downto 0); -- cast44:output -> Avalon_ST_Source_data_0:input
	signal clock_0_clock_output_reset                                 : std_logic;                     -- Clock_0:aclr_out -> [Decoder1:aclr, Decoder:aclr, Delay1:aclr, Delay2:aclr, Delay3:aclr, Delay:aclr, Test_Pattern_Generator_CTRL_PAK_TRANSLATE_0:aclr, Test_Pattern_Generator_DATA_GENERATE_0:aclr, Test_Pattern_Generator_MAIN_CTRL_0:aclr]
	signal clock_0_clock_output_clk                                   : std_logic;                     -- Clock_0:clock_out -> [Decoder1:clock, Decoder:clock, Delay1:clock, Delay2:clock, Delay3:clock, Delay:clock, Test_Pattern_Generator_CTRL_PAK_TRANSLATE_0:Clock, Test_Pattern_Generator_DATA_GENERATE_0:Clock, Test_Pattern_Generator_MAIN_CTRL_0:Clock]

begin

	clock_0 : component alt_dspbuilder_clock_GNF343OQUJ
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr_n    => aclr                        --             .reset_n
		);

	avalon_mm_slave_address_0 : component alt_dspbuilder_port_GN6TDLHAW6
		port map (
			input  => Avalon_MM_Slave_address,               --  input.wire
			output => avalon_mm_slave_address_0_output_wire  -- output.wire
		);

	test_pattern_generator_data_generate_0 : component Test_Pattern_Generator_GN_Test_Pattern_Generator_DATA_GENERATE
		port map (
			Clock    => clock_0_clock_output_clk,                             --    Clock.clk
			aclr     => clock_0_clock_output_reset,                           --         .reset
			counter  => test_pattern_generator_main_ctrl_0_counter_1_wire,    --  counter.wire
			col      => delay2_output_wire,                                   --      col.wire
			colorbar => test_pattern_generator_data_generate_0_colorbar_wire, -- colorbar.wire
			data_en  => test_pattern_generator_main_ctrl_0_data_en_wire,      --  data_en.wire
			ctrl_en  => test_pattern_generator_main_ctrl_0_ctrl_en_wire       --  ctrl_en.wire
		);

	avalon_st_source_valid_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => logical_bit_operator2_result_wire, --  input.wire
			output => Avalon_ST_Source_valid             -- output.wire
		);

	avalon_mm_slave_writedata_0 : component alt_dspbuilder_port_GNEPKLLZKY
		port map (
			input  => Avalon_MM_Slave_writedata,               --  input.wire
			output => avalon_mm_slave_writedata_0_output_wire  -- output.wire
		);

	test_pattern_generator_ctrl_pak_translate_0 : component Test_Pattern_Generator_GN_Test_Pattern_Generator_CTRL_PAK_TRANSLATE
		port map (
			ctrl_pak2 => test_pattern_generator_ctrl_pak_translate_0_ctrl_pak2_wire, -- ctrl_pak2.wire
			dil       => constant3_output_wire,                                      --       dil.wire
			col       => delay2_output_wire,                                         --       col.wire
			Clock     => clock_0_clock_output_clk,                                   --     Clock.clk
			aclr      => clock_0_clock_output_reset,                                 --          .reset
			ctrl_pak1 => test_pattern_generator_ctrl_pak_translate_0_ctrl_pak1_wire, -- ctrl_pak1.wire
			ctrl_pak3 => test_pattern_generator_ctrl_pak_translate_0_ctrl_pak3_wire, -- ctrl_pak3.wire
			row       => delay3_output_wire                                          --       row.wire
		);

	avalon_st_source_endofpacket_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => test_pattern_generator_main_ctrl_0_eop_wire, --  input.wire
			output => Avalon_ST_Source_endofpacket                 -- output.wire
		);

	avalon_st_source_startofpacket_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => test_pattern_generator_main_ctrl_0_sop_wire, --  input.wire
			output => Avalon_ST_Source_startofpacket               -- output.wire
		);

	constant3 : component alt_dspbuilder_constant_GNPLBTTHPL
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "0000",
			width      => 4
		)
		port map (
			output => constant3_output_wire  -- output.wire
		);

	delay : component alt_dspbuilder_delay_GNPJ4Y7BVC
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "00000000000000000000000000100000",
			width      => 32
		)
		port map (
			input  => avalon_mm_slave_writedata_0_output_wire, --      input.wire
			clock  => clock_0_clock_output_clk,                -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,              --           .reset
			output => delay_output_wire,                       --     output.wire
			sclr   => delaysclrgnd_output_wire,                --       sclr.wire
			ena    => logical_bit_operator_result_wire         --        ena.wire
		);

	delaysclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delaysclrgnd_output_wire  -- output.wire
		);

	avalon_mm_slave_write_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => Avalon_MM_Slave_write,               --  input.wire
			output => avalon_mm_slave_write_0_output_wire  -- output.wire
		);

	logical_bit_operator2 : component alt_dspbuilder_logical_bit_op_GNUQ2R64DV
		generic map (
			LogicalOp     => "AltOR",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator2_result_wire,               -- result.wire
			data0  => test_pattern_generator_main_ctrl_0_ctrl_en_wire, --  data0.wire
			data1  => test_pattern_generator_main_ctrl_0_data_en_wire  --  data1.wire
		);

	avalon_st_source_data_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => cast44_output_wire,    --  input.wire
			output => Avalon_ST_Source_data  -- output.wire
		);

	logical_bit_operator1 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator1_result_wire,   -- result.wire
			data0  => avalon_mm_slave_write_0_output_wire, --  data0.wire
			data1  => decoder1_dec_wire                    --  data1.wire
		);

	decoder1 : component alt_dspbuilder_decoder_GNEQGKKPXW
		generic map (
			decode   => "10",
			pipeline => 1,
			width    => 2
		)
		port map (
			clock => clock_0_clock_output_clk,              -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset,            --           .reset
			data  => avalon_mm_slave_address_0_output_wire, --       data.wire
			dec   => decoder1_dec_wire,                     --        dec.wire
			sclr  => decoder1sclrgnd_output_wire,           --       sclr.wire
			ena   => decoder1enavcc_output_wire             --        ena.wire
		);

	decoder1sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => decoder1sclrgnd_output_wire  -- output.wire
		);

	decoder1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => decoder1enavcc_output_wire  -- output.wire
		);

	logical_bit_operator : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator_result_wire,    -- result.wire
			data0  => decoder_dec_wire,                    --  data0.wire
			data1  => avalon_mm_slave_write_0_output_wire  --  data1.wire
		);

	test_pattern_generator_main_ctrl_0 : component Test_Pattern_Generator_GN_Test_Pattern_Generator_MAIN_CTRL
		port map (
			eop       => test_pattern_generator_main_ctrl_0_eop_wire,                --       eop.wire
			counter_1 => test_pattern_generator_main_ctrl_0_counter_1_wire,          -- counter_1.wire
			colorbar  => test_pattern_generator_data_generate_0_colorbar_wire,       --  colorbar.wire
			data      => test_pattern_generator_main_ctrl_0_data_wire,               --      data.wire
			col       => delay2_output_wire,                                         --       col.wire
			ctrl_pak3 => test_pattern_generator_ctrl_pak_translate_0_ctrl_pak3_wire, -- ctrl_pak3.wire
			ctrl_pak2 => test_pattern_generator_ctrl_pak_translate_0_ctrl_pak2_wire, -- ctrl_pak2.wire
			data_en   => test_pattern_generator_main_ctrl_0_data_en_wire,            --   data_en.wire
			ctrl_en   => test_pattern_generator_main_ctrl_0_ctrl_en_wire,            --   ctrl_en.wire
			Clock     => clock_0_clock_output_clk,                                   --     Clock.clk
			aclr      => clock_0_clock_output_reset,                                 --          .reset
			row       => delay3_output_wire,                                         --       row.wire
			ctrl_pak1 => test_pattern_generator_ctrl_pak_translate_0_ctrl_pak1_wire, -- ctrl_pak1.wire
			check_en  => test_pattern_generator_main_ctrl_0_check_en_wire,           --  check_en.wire
			sop       => test_pattern_generator_main_ctrl_0_sop_wire,                --       sop.wire
			ready     => avalon_st_source_ready_0_output_wire                        --     ready.wire
		);

	delay3 : component alt_dspbuilder_delay_GNPJ4Y7BVC
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "00000000000000000000000000100000",
			width      => 32
		)
		port map (
			input  => delay1_output_wire,                               --      input.wire
			clock  => clock_0_clock_output_clk,                         -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,                       --           .reset
			output => delay3_output_wire,                               --     output.wire
			sclr   => delay3sclrgnd_output_wire,                        --       sclr.wire
			ena    => test_pattern_generator_main_ctrl_0_check_en_wire  --        ena.wire
		);

	delay3sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay3sclrgnd_output_wire  -- output.wire
		);

	delay1 : component alt_dspbuilder_delay_GNPJ4Y7BVC
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "00000000000000000000000000100000",
			width      => 32
		)
		port map (
			input  => avalon_mm_slave_writedata_0_output_wire, --      input.wire
			clock  => clock_0_clock_output_clk,                -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,              --           .reset
			output => delay1_output_wire,                      --     output.wire
			sclr   => delay1sclrgnd_output_wire,               --       sclr.wire
			ena    => logical_bit_operator1_result_wire        --        ena.wire
		);

	delay1sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay1sclrgnd_output_wire  -- output.wire
		);

	delay2 : component alt_dspbuilder_delay_GNPJ4Y7BVC
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 1,
			BitPattern => "00000000000000000000000000100000",
			width      => 32
		)
		port map (
			input  => delay_output_wire,                                --      input.wire
			clock  => clock_0_clock_output_clk,                         -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,                       --           .reset
			output => delay2_output_wire,                               --     output.wire
			sclr   => delay2sclrgnd_output_wire,                        --       sclr.wire
			ena    => test_pattern_generator_main_ctrl_0_check_en_wire  --        ena.wire
		);

	delay2sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay2sclrgnd_output_wire  -- output.wire
		);

	avalon_st_source_ready_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => Avalon_ST_Source_ready,               --  input.wire
			output => avalon_st_source_ready_0_output_wire  -- output.wire
		);

	decoder : component alt_dspbuilder_decoder_GNM4LOIHXZ
		generic map (
			decode   => "01",
			pipeline => 1,
			width    => 2
		)
		port map (
			clock => clock_0_clock_output_clk,              -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset,            --           .reset
			data  => avalon_mm_slave_address_0_output_wire, --       data.wire
			dec   => decoder_dec_wire,                      --        dec.wire
			sclr  => decodersclrgnd_output_wire,            --       sclr.wire
			ena   => decoderenavcc_output_wire              --        ena.wire
		);

	decodersclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => decodersclrgnd_output_wire  -- output.wire
		);

	decoderenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => decoderenavcc_output_wire  -- output.wire
		);

	cast44 : component alt_dspbuilder_cast_GN5EYRLJQW
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => test_pattern_generator_main_ctrl_0_data_wire, --  input.wire
			output => cast44_output_wire                            -- output.wire
		);

end architecture rtl; -- of Test_Pattern_Generator_GN
