-- Test_Pattern_Generator_GN_Test_Pattern_Generator_DATA_GENERATE.vhd

-- Generated using ACDS version 13.1 162 at 2015.02.11.10:36:05

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Test_Pattern_Generator_GN_Test_Pattern_Generator_DATA_GENERATE is
	port (
		data_en  : in  std_logic                     := '0';             --  data_en.wire
		Clock    : in  std_logic                     := '0';             --    Clock.clk
		aclr     : in  std_logic                     := '0';             --         .reset
		col      : in  std_logic_vector(31 downto 0) := (others => '0'); --      col.wire
		ctrl_en  : in  std_logic                     := '0';             --  ctrl_en.wire
		colorbar : out std_logic_vector(23 downto 0);                    -- colorbar.wire
		counter  : in  std_logic_vector(23 downto 0) := (others => '0')  --  counter.wire
	);
end entity Test_Pattern_Generator_GN_Test_Pattern_Generator_DATA_GENERATE;

architecture rtl of Test_Pattern_Generator_GN_Test_Pattern_Generator_DATA_GENERATE is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_pipelined_adder_GNWEIMU3MK is
		generic (
			width    : natural := 0;
			pipeline : integer := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GNWEIMU3MK;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_port_GNEPKLLZKY is
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNEPKLLZKY;

	component alt_dspbuilder_bus_build_GNI6E4JZ66 is
		generic (
			width : natural := 8
		);
		port (
			output : out std_logic_vector(2 downto 0);        -- wire
			in0    : in  std_logic                    := 'X'; -- wire
			in1    : in  std_logic                    := 'X'; -- wire
			in2    : in  std_logic                    := 'X'  -- wire
		);
	end component alt_dspbuilder_bus_build_GNI6E4JZ66;

	component alt_dspbuilder_divider_GNKAPZN5MO is
		generic (
			Signed   : natural := 0;
			width    : natural := 8;
			pipeline : natural := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			clock     : in  std_logic                          := 'X';             -- clk
			denom     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			numer     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			quotient  : out std_logic_vector(width-1 downto 0);                    -- wire
			remain    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_divider_GNKAPZN5MO;

	component alt_dspbuilder_port_GNOC3SGKQJ is
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNOC3SGKQJ;

	component alt_dspbuilder_if_statement_GNJ7D74ANQ is
		generic (
			use_else_output : natural := 0;
			bwr             : natural := 0;
			use_else_input  : natural := 0;
			signed          : natural := 1;
			HDLTYPE         : string  := "STD_LOGIC_VECTOR";
			if_expression   : string  := "a";
			number_inputs   : integer := 1;
			width           : natural := 8
		);
		port (
			true : out std_logic;                                        -- wire
			a    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			b    : in  std_logic_vector(23 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_if_statement_GNJ7D74ANQ;

	component alt_dspbuilder_constant_GNKT7L5CDY is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNKT7L5CDY;

	component alt_dspbuilder_if_statement_GNIV4UP6ZO is
		generic (
			use_else_output : natural := 0;
			bwr             : natural := 0;
			use_else_input  : natural := 0;
			signed          : natural := 1;
			HDLTYPE         : string  := "STD_LOGIC_VECTOR";
			if_expression   : string  := "a";
			number_inputs   : integer := 1;
			width           : natural := 8
		);
		port (
			true : out std_logic;                                        -- wire
			a    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			b    : in  std_logic_vector(23 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_if_statement_GNIV4UP6ZO;

	component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'; -- wire
			data1  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V;

	component alt_dspbuilder_if_statement_GNMQPB5LUF is
		generic (
			use_else_output : natural := 0;
			bwr             : natural := 0;
			use_else_input  : natural := 0;
			signed          : natural := 1;
			HDLTYPE         : string  := "STD_LOGIC_VECTOR";
			if_expression   : string  := "a";
			number_inputs   : integer := 1;
			width           : natural := 8
		);
		port (
			true : out std_logic;                                        -- wire
			a    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			b    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			c    : in  std_logic_vector(23 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_if_statement_GNMQPB5LUF;

	component alt_dspbuilder_if_statement_GNZR777PB6 is
		generic (
			use_else_output : natural := 0;
			bwr             : natural := 0;
			use_else_input  : natural := 0;
			signed          : natural := 1;
			HDLTYPE         : string  := "STD_LOGIC_VECTOR";
			if_expression   : string  := "a";
			number_inputs   : integer := 1;
			width           : natural := 8
		);
		port (
			true : out std_logic;                                        -- wire
			a    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			b    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			c    : in  std_logic_vector(23 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_if_statement_GNZR777PB6;

	component alt_dspbuilder_constant_GNUWBUDS4L is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNUWBUDS4L;

	component alt_dspbuilder_constant_GNJ2DIDH6N is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNJ2DIDH6N;

	component alt_dspbuilder_logical_bit_op_GNUQ2R64DV is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'; -- wire
			data1  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNUQ2R64DV;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_constant_GNNCFWNIJI is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(15 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNNCFWNIJI;

	component alt_dspbuilder_if_statement_GNWHMBR6GA is
		generic (
			use_else_output : natural := 0;
			bwr             : natural := 0;
			use_else_input  : natural := 0;
			signed          : natural := 1;
			HDLTYPE         : string  := "STD_LOGIC_VECTOR";
			if_expression   : string  := "a";
			number_inputs   : integer := 1;
			width           : natural := 8
		);
		port (
			true : out std_logic;                                        -- wire
			a    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			b    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			c    : in  std_logic_vector(23 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_if_statement_GNWHMBR6GA;

	component alt_dspbuilder_single_pulse_GN2XGKTRR3 is
		generic (
			delay         : positive := 1;
			signal_type   : string   := "Impulse";
			impulse_width : positive := 1
		);
		port (
			aclr   : in  std_logic := 'X'; -- clk
			clock  : in  std_logic := 'X'; -- clk
			ena    : in  std_logic := 'X'; -- wire
			result : out std_logic;        -- wire
			sclr   : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_single_pulse_GN2XGKTRR3;

	component StateMachineEditor1 is
		port (
			clock      : in  std_logic                     := 'X';             -- clk
			col_select : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- wire
			data       : out std_logic_vector(23 downto 0);                    -- wire
			data_en    : in  std_logic                     := 'X';             -- wire
			reset      : in  std_logic                     := 'X'              -- wire
		);
	end component StateMachineEditor1;

	component alt_dspbuilder_counter_GNZKRIGTBB is
		generic (
			use_usr_aclr : string  := "false";
			use_ena      : string  := "false";
			use_cin      : string  := "false";
			use_sset     : string  := "false";
			ndirection   : natural := 1;
			svalue       : string  := "0";
			use_sload    : string  := "false";
			use_sclr     : string  := "false";
			use_cout     : string  := "false";
			modulus      : integer := 256;
			use_cnt_ena  : string  := "false";
			width        : natural := 8;
			use_aset     : string  := "false";
			use_aload    : string  := "false";
			avalue       : string  := "0"
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			aload     : in  std_logic                          := 'X';             -- wire
			aset      : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cnt_ena   : in  std_logic                          := 'X';             -- wire
			cout      : out std_logic;                                             -- wire
			data      : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			direction : in  std_logic                          := 'X';             -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			q         : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr      : in  std_logic                          := 'X';             -- wire
			sload     : in  std_logic                          := 'X';             -- wire
			sset      : in  std_logic                          := 'X';             -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_counter_GNZKRIGTBB;

	component alt_dspbuilder_multiplier_GNEIWYOKUR is
		generic (
			DEDICATED_MULTIPLIER_CIRCUITRY : string  := "AUTO";
			Signed                         : natural := 0;
			OutputMsb                      : integer := 8;
			aWidth                         : natural := 8;
			bWidth                         : natural := 8;
			OutputLsb                      : integer := 0;
			pipeline                       : integer := 0
		);
		port (
			aclr      : in  std_logic                                          := 'X';             -- clk
			clock     : in  std_logic                                          := 'X';             -- clk
			dataa     : in  std_logic_vector(aWidth-1 downto 0)                := (others => 'X'); -- wire
			datab     : in  std_logic_vector(bWidth-1 downto 0)                := (others => 'X'); -- wire
			ena       : in  std_logic                                          := 'X';             -- wire
			result    : out std_logic_vector(OutputMsb-OutputLsb+1-1 downto 0);                    -- wire
			user_aclr : in  std_logic                                          := 'X'              -- wire
		);
	end component alt_dspbuilder_multiplier_GNEIWYOKUR;

	component alt_dspbuilder_cast_GN7PRGDOVA is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN7PRGDOVA;

	component alt_dspbuilder_cast_GNCPEUNC4M is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNCPEUNC4M;

	component alt_dspbuilder_cast_GNKIWLRTQI is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(47 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNKIWLRTQI;

	component alt_dspbuilder_cast_GNLHWQIRQK is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(2 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(2 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNLHWQIRQK;

	signal pipelined_adder3user_aclrgnd_output_wire : std_logic;                     -- Pipelined_Adder3user_aclrGND:output -> Pipelined_Adder3:user_aclr
	signal pipelined_adder3enavcc_output_wire       : std_logic;                     -- Pipelined_Adder3enaVCC:output -> Pipelined_Adder3:ena
	signal divideruser_aclrgnd_output_wire          : std_logic;                     -- Divideruser_aclrGND:output -> Divider:user_aclr
	signal dividerenavcc_output_wire                : std_logic;                     -- DividerenaVCC:output -> Divider:ena
	signal single_pulse1sclrgnd_output_wire         : std_logic;                     -- Single_Pulse1sclrGND:output -> Single_Pulse1:sclr
	signal single_pulse1enavcc_output_wire          : std_logic;                     -- Single_Pulse1enaVCC:output -> Single_Pulse1:ena
	signal multiplieruser_aclrgnd_output_wire       : std_logic;                     -- Multiplieruser_aclrGND:output -> Multiplier:user_aclr
	signal multiplierenavcc_output_wire             : std_logic;                     -- MultiplierenaVCC:output -> Multiplier:ena
	signal constant9_output_wire                    : std_logic_vector(23 downto 0); -- Constant9:output -> Counter1:data
	signal constant8_output_wire                    : std_logic_vector(23 downto 0); -- Constant8:output -> Divider:denom
	signal counter1_q_wire                          : std_logic_vector(23 downto 0); -- Counter1:q -> [If_Statement1:a, If_Statement2:a, If_Statement3:a, If_Statement:a]
	signal divider_quotient_wire                    : std_logic_vector(23 downto 0); -- Divider:quotient -> [If_Statement1:b, If_Statement:b, Multiplier:dataa]
	signal if_statement_true_wire                   : std_logic;                     -- If_Statement:true -> Bus_Builder:in0
	signal if_statement1_true_wire                  : std_logic;                     -- If_Statement1:true -> Bus_Builder:in1
	signal if_statement2_true_wire                  : std_logic;                     -- If_Statement2:true -> Bus_Builder:in2
	signal counter_0_output_wire                    : std_logic_vector(23 downto 0); -- counter_0:output -> If_Statement5:a
	signal if_statement3_true_wire                  : std_logic;                     -- If_Statement3:true -> Logical_Bit_Operator12:data0
	signal data_en_0_output_wire                    : std_logic;                     -- data_en_0:output -> [Logical_Bit_Operator12:data1, Logical_Bit_Operator8:data0, State_Machine_Editor1:data_en]
	signal ctrl_en_0_output_wire                    : std_logic;                     -- ctrl_en_0:output -> Logical_Bit_Operator7:data0
	signal logical_bit_operator12_result_wire       : std_logic;                     -- Logical_Bit_Operator12:result -> Logical_Bit_Operator7:data1
	signal logical_bit_operator7_result_wire        : std_logic;                     -- Logical_Bit_Operator7:result -> Counter1:sload
	signal if_statement5_true_wire                  : std_logic;                     -- If_Statement5:true -> Logical_Bit_Operator8:data1
	signal logical_bit_operator8_result_wire        : std_logic;                     -- Logical_Bit_Operator8:result -> Counter1:cnt_ena
	signal constant6_output_wire                    : std_logic_vector(23 downto 0); -- Constant6:output -> Multiplier:datab
	signal constant13_output_wire                   : std_logic_vector(23 downto 0); -- Constant13:output -> Pipelined_Adder3:datab
	signal pipelined_adder3_result_wire             : std_logic_vector(23 downto 0); -- Pipelined_Adder3:result -> If_Statement2:c
	signal single_pulse1_result_wire                : std_logic;                     -- Single_Pulse1:result -> State_Machine_Editor1:reset
	signal state_machine_editor1_data_wire          : std_logic_vector(23 downto 0); -- State_Machine_Editor1:data -> colorbar_0:input
	signal col_0_output_wire                        : std_logic_vector(31 downto 0); -- col_0:output -> [cast0:input, cast1:input, cast2:input, cast6:input]
	signal cast0_output_wire                        : std_logic_vector(23 downto 0); -- cast0:output -> Divider:numer
	signal cast1_output_wire                        : std_logic_vector(23 downto 0); -- cast1:output -> If_Statement:c
	signal cast2_output_wire                        : std_logic_vector(23 downto 0); -- cast2:output -> If_Statement3:b
	signal constant11_output_wire                   : std_logic_vector(15 downto 0); -- Constant11:output -> cast3:input
	signal cast3_output_wire                        : std_logic_vector(23 downto 0); -- cast3:output -> If_Statement5:b
	signal multiplier_result_wire                   : std_logic_vector(47 downto 0); -- Multiplier:result -> [cast4:input, cast5:input]
	signal cast4_output_wire                        : std_logic_vector(23 downto 0); -- cast4:output -> If_Statement1:c
	signal cast5_output_wire                        : std_logic_vector(23 downto 0); -- cast5:output -> If_Statement2:b
	signal cast6_output_wire                        : std_logic_vector(23 downto 0); -- cast6:output -> Pipelined_Adder3:dataa
	signal bus_builder_output_wire                  : std_logic_vector(2 downto 0);  -- Bus_Builder:output -> cast7:input
	signal cast7_output_wire                        : std_logic_vector(2 downto 0);  -- cast7:output -> State_Machine_Editor1:col_select
	signal clock_0_clock_output_reset               : std_logic;                     -- Clock_0:aclr_out -> [Counter1:aclr, Divider:aclr, Multiplier:aclr, Pipelined_Adder3:aclr, Single_Pulse1:aclr]
	signal clock_0_clock_output_clk                 : std_logic;                     -- Clock_0:clock_out -> [Counter1:clock, Divider:clock, Multiplier:clock, Pipelined_Adder3:clock, Single_Pulse1:clock, State_Machine_Editor1:clock]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	pipelined_adder3 : component alt_dspbuilder_pipelined_adder_GNWEIMU3MK
		generic map (
			width    => 24,
			pipeline => 2
		)
		port map (
			clock     => clock_0_clock_output_clk,                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,               --           .reset
			dataa     => cast6_output_wire,                        --      dataa.wire
			datab     => constant13_output_wire,                   --      datab.wire
			result    => pipelined_adder3_result_wire,             --     result.wire
			user_aclr => pipelined_adder3user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder3enavcc_output_wire        --        ena.wire
		);

	pipelined_adder3user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder3user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder3enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder3enavcc_output_wire  -- output.wire
		);

	col_0 : component alt_dspbuilder_port_GNEPKLLZKY
		port map (
			input  => col,               --  input.wire
			output => col_0_output_wire  -- output.wire
		);

	bus_builder : component alt_dspbuilder_bus_build_GNI6E4JZ66
		generic map (
			width => 3
		)
		port map (
			output => bus_builder_output_wire, -- output.wire
			in0    => if_statement_true_wire,  --    in0.wire
			in1    => if_statement1_true_wire, --    in1.wire
			in2    => if_statement2_true_wire  --    in2.wire
		);

	divider : component alt_dspbuilder_divider_GNKAPZN5MO
		generic map (
			Signed   => 0,
			width    => 24,
			pipeline => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,        -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,      --           .reset
			numer     => cast0_output_wire,               --      numer.wire
			denom     => constant8_output_wire,           --      denom.wire
			quotient  => divider_quotient_wire,           --   quotient.wire
			remain    => open,                            --     remain.wire
			user_aclr => divideruser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => dividerenavcc_output_wire        --        ena.wire
		);

	divideruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => divideruser_aclrgnd_output_wire  -- output.wire
		);

	dividerenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => dividerenavcc_output_wire  -- output.wire
		);

	colorbar_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => state_machine_editor1_data_wire, --  input.wire
			output => colorbar                         -- output.wire
		);

	if_statement5 : component alt_dspbuilder_if_statement_GNJ7D74ANQ
		generic map (
			use_else_output => 0,
			bwr             => 0,
			use_else_input  => 0,
			signed          => 0,
			HDLTYPE         => "STD_LOGIC_VECTOR",
			if_expression   => "a>b",
			number_inputs   => 2,
			width           => 24
		)
		port map (
			true => if_statement5_true_wire, -- true.wire
			a    => counter_0_output_wire,   --    a.wire
			b    => cast3_output_wire        --    b.wire
		);

	counter_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => counter,               --  input.wire
			output => counter_0_output_wire  -- output.wire
		);

	constant6 : component alt_dspbuilder_constant_GNKT7L5CDY
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "000000000000000000000010",
			width      => 24
		)
		port map (
			output => constant6_output_wire  -- output.wire
		);

	if_statement3 : component alt_dspbuilder_if_statement_GNIV4UP6ZO
		generic map (
			use_else_output => 0,
			bwr             => 0,
			use_else_input  => 0,
			signed          => 0,
			HDLTYPE         => "STD_LOGIC_VECTOR",
			if_expression   => "a=b",
			number_inputs   => 2,
			width           => 24
		)
		port map (
			true => if_statement3_true_wire, -- true.wire
			a    => counter1_q_wire,         --    a.wire
			b    => cast2_output_wire        --    b.wire
		);

	logical_bit_operator12 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator12_result_wire, -- result.wire
			data0  => if_statement3_true_wire,            --  data0.wire
			data1  => data_en_0_output_wire               --  data1.wire
		);

	if_statement2 : component alt_dspbuilder_if_statement_GNMQPB5LUF
		generic map (
			use_else_output => 0,
			bwr             => 0,
			use_else_input  => 0,
			signed          => 0,
			HDLTYPE         => "STD_LOGIC_VECTOR",
			if_expression   => "((a>b) or (a=b)) and ((a<c) or (a=c))",
			number_inputs   => 3,
			width           => 24
		)
		port map (
			true => if_statement2_true_wire,      -- true.wire
			a    => counter1_q_wire,              --    a.wire
			b    => cast5_output_wire,            --    b.wire
			c    => pipelined_adder3_result_wire  --    c.wire
		);

	if_statement1 : component alt_dspbuilder_if_statement_GNZR777PB6
		generic map (
			use_else_output => 0,
			bwr             => 0,
			use_else_input  => 0,
			signed          => 0,
			HDLTYPE         => "STD_LOGIC_VECTOR",
			if_expression   => "((a>b) or (a=b)) and (a<c)",
			number_inputs   => 3,
			width           => 24
		)
		port map (
			true => if_statement1_true_wire, -- true.wire
			a    => counter1_q_wire,         --    a.wire
			b    => divider_quotient_wire,   --    b.wire
			c    => cast4_output_wire        --    c.wire
		);

	constant8 : component alt_dspbuilder_constant_GNUWBUDS4L
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "000000000000000000000011",
			width      => 24
		)
		port map (
			output => constant8_output_wire  -- output.wire
		);

	constant9 : component alt_dspbuilder_constant_GNJ2DIDH6N
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "000000000000000000000001",
			width      => 24
		)
		port map (
			output => constant9_output_wire  -- output.wire
		);

	logical_bit_operator7 : component alt_dspbuilder_logical_bit_op_GNUQ2R64DV
		generic map (
			LogicalOp     => "AltOR",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator7_result_wire,  -- result.wire
			data0  => ctrl_en_0_output_wire,              --  data0.wire
			data1  => logical_bit_operator12_result_wire  --  data1.wire
		);

	ctrl_en_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => ctrl_en,               --  input.wire
			output => ctrl_en_0_output_wire  -- output.wire
		);

	constant11 : component alt_dspbuilder_constant_GNNCFWNIJI
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "0000000000000100",
			width      => 16
		)
		port map (
			output => constant11_output_wire  -- output.wire
		);

	if_statement : component alt_dspbuilder_if_statement_GNWHMBR6GA
		generic map (
			use_else_output => 0,
			bwr             => 0,
			use_else_input  => 0,
			signed          => 0,
			HDLTYPE         => "STD_LOGIC_VECTOR",
			if_expression   => "((a>zero) and (a<b)) or (a=c)",
			number_inputs   => 3,
			width           => 24
		)
		port map (
			true => if_statement_true_wire, -- true.wire
			a    => counter1_q_wire,        --    a.wire
			b    => divider_quotient_wire,  --    b.wire
			c    => cast1_output_wire       --    c.wire
		);

	data_en_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => data_en,               --  input.wire
			output => data_en_0_output_wire  -- output.wire
		);

	constant13 : component alt_dspbuilder_constant_GNJ2DIDH6N
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "000000000000000000000001",
			width      => 24
		)
		port map (
			output => constant13_output_wire  -- output.wire
		);

	logical_bit_operator8 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator8_result_wire, -- result.wire
			data0  => data_en_0_output_wire,             --  data0.wire
			data1  => if_statement5_true_wire            --  data1.wire
		);

	single_pulse1 : component alt_dspbuilder_single_pulse_GN2XGKTRR3
		generic map (
			delay         => 1,
			signal_type   => "Step Down",
			impulse_width => 1
		)
		port map (
			clock  => clock_0_clock_output_clk,         -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,       --           .reset
			result => single_pulse1_result_wire,        --     result.wire
			sclr   => single_pulse1sclrgnd_output_wire, --       sclr.wire
			ena    => single_pulse1enavcc_output_wire   --        ena.wire
		);

	single_pulse1sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => single_pulse1sclrgnd_output_wire  -- output.wire
		);

	single_pulse1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => single_pulse1enavcc_output_wire  -- output.wire
		);

	state_machine_editor1 : component StateMachineEditor1
		port map (
			clock      => clock_0_clock_output_clk,        --      clock.clk
			reset      => single_pulse1_result_wire,       --      reset.wire
			col_select => cast7_output_wire,               -- col_select.wire
			data_en    => data_en_0_output_wire,           --    data_en.wire
			data       => state_machine_editor1_data_wire  --       data.wire
		);

	counter1 : component alt_dspbuilder_counter_GNZKRIGTBB
		generic map (
			use_usr_aclr => "false",
			use_ena      => "false",
			use_cin      => "false",
			use_sset     => "false",
			ndirection   => 1,
			svalue       => "1",
			use_sload    => "true",
			use_sclr     => "false",
			use_cout     => "false",
			modulus      => 65536,
			use_cnt_ena  => "true",
			width        => 24,
			use_aset     => "false",
			use_aload    => "false",
			avalue       => "0"
		)
		port map (
			clock   => clock_0_clock_output_clk,          -- clock_aclr.clk
			aclr    => clock_0_clock_output_reset,        --           .reset
			data    => constant9_output_wire,             --       data.wire
			cnt_ena => logical_bit_operator8_result_wire, --    cnt_ena.wire
			sload   => logical_bit_operator7_result_wire, --      sload.wire
			q       => counter1_q_wire,                   --          q.wire
			cout    => open                               --       cout.wire
		);

	multiplier : component alt_dspbuilder_multiplier_GNEIWYOKUR
		generic map (
			DEDICATED_MULTIPLIER_CIRCUITRY => "YES",
			Signed                         => 0,
			OutputMsb                      => 47,
			aWidth                         => 24,
			bWidth                         => 24,
			OutputLsb                      => 0,
			pipeline                       => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,           -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,         --           .reset
			dataa     => divider_quotient_wire,              --      dataa.wire
			datab     => constant6_output_wire,              --      datab.wire
			result    => multiplier_result_wire,             --     result.wire
			user_aclr => multiplieruser_aclrgnd_output_wire, --  user_aclr.wire
			ena       => multiplierenavcc_output_wire        --        ena.wire
		);

	multiplieruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplieruser_aclrgnd_output_wire  -- output.wire
		);

	multiplierenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplierenavcc_output_wire  -- output.wire
		);

	cast0 : component alt_dspbuilder_cast_GN7PRGDOVA
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => col_0_output_wire, --  input.wire
			output => cast0_output_wire  -- output.wire
		);

	cast1 : component alt_dspbuilder_cast_GN7PRGDOVA
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => col_0_output_wire, --  input.wire
			output => cast1_output_wire  -- output.wire
		);

	cast2 : component alt_dspbuilder_cast_GN7PRGDOVA
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => col_0_output_wire, --  input.wire
			output => cast2_output_wire  -- output.wire
		);

	cast3 : component alt_dspbuilder_cast_GNCPEUNC4M
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant11_output_wire, --  input.wire
			output => cast3_output_wire       -- output.wire
		);

	cast4 : component alt_dspbuilder_cast_GNKIWLRTQI
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier_result_wire, --  input.wire
			output => cast4_output_wire       -- output.wire
		);

	cast5 : component alt_dspbuilder_cast_GNKIWLRTQI
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier_result_wire, --  input.wire
			output => cast5_output_wire       -- output.wire
		);

	cast6 : component alt_dspbuilder_cast_GN7PRGDOVA
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => col_0_output_wire, --  input.wire
			output => cast6_output_wire  -- output.wire
		);

	cast7 : component alt_dspbuilder_cast_GNLHWQIRQK
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => bus_builder_output_wire, --  input.wire
			output => cast7_output_wire        -- output.wire
		);

end architecture rtl; -- of Test_Pattern_Generator_GN_Test_Pattern_Generator_DATA_GENERATE
