-- Copyright (C) 1991-2013 Altera Corporation
-- Your use of Altera Corporation's design tools, logic functions 
-- and other software and tools, and its AMPP partner logic 
-- functions, and any output files from any of the foregoing 
-- (including device programming or simulation files), and any 
-- associated documentation or information are expressly subject 
-- to the terms and conditions of the Altera Program License 
-- Subscription Agreement, Altera MegaCore Function License 
-- Agreement, or other applicable license agreement, including, 
-- without limitation, that your use is for the sole purpose of 
-- programming logic devices manufactured by Altera and sold by 
-- Altera or its authorized distributors.  Please refer to the 
-- applicable agreement for further details.

-- Generated by Quartus II Version 13.1.0 Build 162 10/23/2013 SJ Full Version
-- Created on Wed Feb 11 10:17:50 2015

LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY StateMachineEditor IS
    PORT (
        clock : IN STD_LOGIC;
        reset : IN STD_LOGIC := '0';
        ready : IN STD_LOGIC := '0';
        counter : IN STD_LOGIC_VECTOR(23 DOWNTO 0) := "000000000000000000000000";
        data_end : IN STD_LOGIC := '0';
        state : OUT STD_LOGIC_VECTOR(2 DOWNTO 0)
    );
END StateMachineEditor;

ARCHITECTURE BEHAVIOR OF StateMachineEditor IS
    TYPE type_fstate IS (CTRL,DATA,IDLE);
    SIGNAL fstate : type_fstate;
    SIGNAL reg_fstate : type_fstate;
BEGIN
    PROCESS (clock,reg_fstate)
    BEGIN
        IF (clock='1' AND clock'event) THEN
            fstate <= reg_fstate;
        END IF;
    END PROCESS;

    PROCESS (fstate,reset,ready,counter,data_end)
    BEGIN
        IF (reset='1') THEN
            reg_fstate <= IDLE;
            state <= "000";
        ELSE
            state <= "000";
            CASE fstate IS
                WHEN CTRL =>
                    IF (((ready = '0') OR (counter(23 DOWNTO 0) = "000000000000000000000011"))) THEN
                        reg_fstate <= IDLE;
                    ELSIF (((ready = '1') AND (counter(23 DOWNTO 0) < "000000000000000000000011"))) THEN
                        reg_fstate <= CTRL;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= CTRL;
                    END IF;

                    state <= "001";
                WHEN DATA =>
                    IF (((ready = '0') OR ((ready = '1') AND (data_end = '1')))) THEN
                        reg_fstate <= IDLE;
                    ELSIF (((ready = '1') AND (data_end = '0'))) THEN
                        reg_fstate <= DATA;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= DATA;
                    END IF;

                    state <= "010";
                WHEN IDLE =>
                    IF (((ready = '1') AND (counter(23 DOWNTO 0) > "000000000000000000000011"))) THEN
                        reg_fstate <= DATA;
                    ELSIF (((ready = '1') AND (counter(23 DOWNTO 0) <= "000000000000000000000011"))) THEN
                        reg_fstate <= CTRL;
                    ELSIF ((ready = '0')) THEN
                        reg_fstate <= IDLE;
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        reg_fstate <= IDLE;
                    END IF;

                    IF ((counter(23 DOWNTO 0) /= "000000000000000000000000")) THEN
                        state <= "000";
                    ELSIF ((counter(23 DOWNTO 0) = "000000000000000000000000")) THEN
                        state <= "100";
                    -- Inserting 'else' block to prevent latch inference
                    ELSE
                        state <= "000";
                    END IF;
                WHEN OTHERS => 
                    state <= "XXX";
                    report "Reach undefined state";
            END CASE;
        END IF;
    END PROCESS;
END BEHAVIOR;
