-- Test_Pattern_Generator_GN_Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT.vhd

-- Generated using ACDS version 13.1 162 at 2015.02.11.10:36:06

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Test_Pattern_Generator_GN_Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT is
	port (
		eop       : out std_logic;                                        --       eop.wire
		data_en   : in  std_logic                     := '0';             --   data_en.wire
		ctrl_pak3 : in  std_logic_vector(23 downto 0) := (others => '0'); -- ctrl_pak3.wire
		ctrl_pak1 : in  std_logic_vector(23 downto 0) := (others => '0'); -- ctrl_pak1.wire
		ctrl_en   : in  std_logic                     := '0';             --   ctrl_en.wire
		sop       : out std_logic;                                        --       sop.wire
		data      : out std_logic_vector(24 downto 0);                    --      data.wire
		ctrl_pak2 : in  std_logic_vector(23 downto 0) := (others => '0'); -- ctrl_pak2.wire
		pixel_num : in  std_logic_vector(47 downto 0) := (others => '0'); -- pixel_num.wire
		colorbar  : in  std_logic_vector(23 downto 0) := (others => '0'); --  colorbar.wire
		counter   : in  std_logic_vector(23 downto 0) := (others => '0'); --   counter.wire
		Clock     : in  std_logic                     := '0';             --     Clock.clk
		aclr      : in  std_logic                     := '0'              --          .reset
	);
end entity Test_Pattern_Generator_GN_Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT;

architecture rtl of Test_Pattern_Generator_GN_Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_cast_GN33BXJAZX is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(1 downto 0)                      -- wire
		);
	end component alt_dspbuilder_cast_GN33BXJAZX;

	component alt_dspbuilder_pipelined_adder_GNTWZRTG4I is
		generic (
			width    : natural := 0;
			pipeline : integer := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GNTWZRTG4I;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_case_statement_GNWMX2GCN2 is
		generic (
			number_outputs : integer := 8;
			hasDefault     : natural := 0;
			pipeline       : natural := 0;
			width          : integer := 8
		);
		port (
			clock : in  std_logic                     := 'X';             -- clk
			aclr  : in  std_logic                     := 'X';             -- reset
			input : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			r0    : out std_logic;                                        -- wire
			r1    : out std_logic                                         -- wire
		);
	end component alt_dspbuilder_case_statement_GNWMX2GCN2;

	component alt_dspbuilder_case_statement_GNFTM45DFU is
		generic (
			number_outputs : integer := 8;
			hasDefault     : natural := 0;
			pipeline       : natural := 0;
			width          : integer := 8
		);
		port (
			clock : in  std_logic                     := 'X';             -- clk
			aclr  : in  std_logic                     := 'X';             -- reset
			input : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			r0    : out std_logic;                                        -- wire
			r1    : out std_logic                                         -- wire
		);
	end component alt_dspbuilder_case_statement_GNFTM45DFU;

	component alt_dspbuilder_multiplexer_GNLGLCKYZ5 is
		generic (
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0;
			width                  : positive := 8;
			pipeline               : natural  := 0;
			number_inputs          : natural  := 4
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			sel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- wire
			result    : out std_logic_vector(23 downto 0);                    -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			in0       : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			in2       : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			in3       : in  std_logic_vector(23 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNLGLCKYZ5;

	component alt_dspbuilder_port_GNEHYJMBQS is
		port (
			input  : in  std_logic_vector(24 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(24 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNEHYJMBQS;

	component alt_dspbuilder_constant_GNNKZSYI73 is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNNKZSYI73;

	component alt_dspbuilder_bus_concat_GN6E6AAQPZ is
		generic (
			widthB : natural := 8;
			widthA : natural := 8
		);
		port (
			a      : in  std_logic_vector(widthA-1 downto 0)        := (others => 'X'); -- wire
			aclr   : in  std_logic                                  := 'X';             -- clk
			b      : in  std_logic_vector(widthB-1 downto 0)        := (others => 'X'); -- wire
			clock  : in  std_logic                                  := 'X';             -- clk
			output : out std_logic_vector(widthA+widthB-1 downto 0)                     -- wire
		);
	end component alt_dspbuilder_bus_concat_GN6E6AAQPZ;

	component alt_dspbuilder_logical_bit_op_GNUQ2R64DV is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'; -- wire
			data1  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNUQ2R64DV;

	component alt_dspbuilder_port_GNOC3SGKQJ is
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNOC3SGKQJ;

	component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'; -- wire
			data1  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V;

	component alt_dspbuilder_constant_GNZEH3JAKA is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNZEH3JAKA;

	component alt_dspbuilder_delay_GNIYBMGPQQ is
		generic (
			ClockPhase : string   := "1";
			delay      : positive := 1;
			use_init   : natural  := 0;
			BitPattern : string   := "00000001";
			width      : positive := 8
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNIYBMGPQQ;

	component alt_dspbuilder_constant_GNLJWFEWBD is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(15 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNLJWFEWBD;

	component alt_dspbuilder_constant_GNQJ63TWA6 is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNQJ63TWA6;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component alt_dspbuilder_if_statement_GNTVBNRAAT is
		generic (
			use_else_output : natural := 0;
			bwr             : natural := 0;
			use_else_input  : natural := 0;
			signed          : natural := 1;
			HDLTYPE         : string  := "STD_LOGIC_VECTOR";
			if_expression   : string  := "a";
			number_inputs   : integer := 1;
			width           : natural := 8
		);
		port (
			true : out std_logic;                                        -- wire
			a    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			b    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			c    : in  std_logic_vector(23 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_if_statement_GNTVBNRAAT;

	component alt_dspbuilder_delay_GNNBTO2F3L is
		generic (
			ClockPhase : string   := "1";
			delay      : positive := 1;
			use_init   : natural  := 0;
			BitPattern : string   := "00000001";
			width      : positive := 8
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNNBTO2F3L;

	component alt_dspbuilder_port_GNUJT4YY5I is
		port (
			input  : in  std_logic_vector(47 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(47 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNUJT4YY5I;

	component alt_dspbuilder_multiplexer_GNHQFFAUXQ is
		generic (
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0;
			width                  : positive := 8;
			pipeline               : natural  := 0;
			number_inputs          : natural  := 4
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			sel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- wire
			result    : out std_logic_vector(24 downto 0);                    -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			in0       : in  std_logic_vector(24 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(24 downto 0) := (others => 'X'); -- wire
			in2       : in  std_logic_vector(24 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GNHQFFAUXQ;

	component alt_dspbuilder_multiplexer_GN6ODCX3D4 is
		generic (
			HDLTYPE                : string   := "STD_LOGIC_VECTOR";
			use_one_hot_select_bus : natural  := 0;
			width                  : positive := 8;
			pipeline               : natural  := 0;
			number_inputs          : natural  := 4
		);
		port (
			clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			sel       : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- wire
			result    : out std_logic_vector(24 downto 0);                    -- wire
			ena       : in  std_logic                     := 'X';             -- wire
			user_aclr : in  std_logic                     := 'X';             -- wire
			in0       : in  std_logic_vector(24 downto 0) := (others => 'X'); -- wire
			in1       : in  std_logic_vector(24 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_multiplexer_GN6ODCX3D4;

	component alt_dspbuilder_delay_GNVJUPFOX3 is
		generic (
			ClockPhase : string   := "1";
			delay      : positive := 1;
			use_init   : natural  := 0;
			BitPattern : string   := "00000001";
			width      : positive := 8
		);
		port (
			aclr   : in  std_logic                          := 'X';             -- clk
			clock  : in  std_logic                          := 'X';             -- clk
			ena    : in  std_logic                          := 'X';             -- wire
			input  : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr   : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_delay_GNVJUPFOX3;

	component alt_dspbuilder_cast_GN3ODVPHOL is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(15 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN3ODVPHOL;

	component alt_dspbuilder_cast_GN46N4UJ5S is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic                    := 'X'; -- wire
			output : out std_logic_vector(0 downto 0)         -- wire
		);
	end component alt_dspbuilder_cast_GN46N4UJ5S;

	component alt_dspbuilder_cast_GNCPEUNC4M is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(15 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNCPEUNC4M;

	component alt_dspbuilder_cast_GNKDE2NVCC is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(24 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNKDE2NVCC;

	component alt_dspbuilder_cast_GNCCZ56SYK is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(24 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNCCZ56SYK;

	component alt_dspbuilder_cast_GNKIWLRTQI is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(47 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNKIWLRTQI;

	signal pipelined_adder2user_aclrgnd_output_wire : std_logic;                     -- Pipelined_Adder2user_aclrGND:output -> Pipelined_Adder2:user_aclr
	signal pipelined_adder2enavcc_output_wire       : std_logic;                     -- Pipelined_Adder2enaVCC:output -> Pipelined_Adder2:ena
	signal multiplexeruser_aclrgnd_output_wire      : std_logic;                     -- Multiplexeruser_aclrGND:output -> Multiplexer:user_aclr
	signal multiplexerenavcc_output_wire            : std_logic;                     -- MultiplexerenaVCC:output -> Multiplexer:ena
	signal delaysclrgnd_output_wire                 : std_logic;                     -- DelaysclrGND:output -> Delay:sclr
	signal delayenavcc_output_wire                  : std_logic;                     -- DelayenaVCC:output -> Delay:ena
	signal delay5sclrgnd_output_wire                : std_logic;                     -- Delay5sclrGND:output -> Delay5:sclr
	signal delay5enavcc_output_wire                 : std_logic;                     -- Delay5enaVCC:output -> Delay5:ena
	signal delay3sclrgnd_output_wire                : std_logic;                     -- Delay3sclrGND:output -> Delay3:sclr
	signal delay3enavcc_output_wire                 : std_logic;                     -- Delay3enaVCC:output -> Delay3:ena
	signal multiplexer1user_aclrgnd_output_wire     : std_logic;                     -- Multiplexer1user_aclrGND:output -> Multiplexer1:user_aclr
	signal multiplexer1enavcc_output_wire           : std_logic;                     -- Multiplexer1enaVCC:output -> Multiplexer1:ena
	signal delay1sclrgnd_output_wire                : std_logic;                     -- Delay1sclrGND:output -> Delay1:sclr
	signal delay1enavcc_output_wire                 : std_logic;                     -- Delay1enaVCC:output -> Delay1:ena
	signal multiplexer2user_aclrgnd_output_wire     : std_logic;                     -- Multiplexer2user_aclrGND:output -> Multiplexer2:user_aclr
	signal multiplexer2enavcc_output_wire           : std_logic;                     -- Multiplexer2enaVCC:output -> Multiplexer2:ena
	signal delay2sclrgnd_output_wire                : std_logic;                     -- Delay2sclrGND:output -> Delay2:sclr
	signal delay2enavcc_output_wire                 : std_logic;                     -- Delay2enaVCC:output -> Delay2:ena
	signal counter_0_output_wire                    : std_logic_vector(23 downto 0); -- counter_0:output -> [Bus_Conversion1:input, If_Statement7:a, cast29:input, cast32:input]
	signal constant1_output_wire                    : std_logic_vector(23 downto 0); -- Constant1:output -> Delay:input
	signal ctrl_pak1_0_output_wire                  : std_logic_vector(23 downto 0); -- ctrl_pak1_0:output -> Delay1:input
	signal ctrl_pak2_0_output_wire                  : std_logic_vector(23 downto 0); -- ctrl_pak2_0:output -> Delay2:input
	signal ctrl_pak3_0_output_wire                  : std_logic_vector(23 downto 0); -- ctrl_pak3_0:output -> Delay3:input
	signal constant7_output_wire                    : std_logic_vector(23 downto 0); -- Constant7:output -> Delay5:input
	signal if_statement7_true_wire                  : std_logic;                     -- If_Statement7:true -> [Logical_Bit_Operator10:data0, Logical_Bit_Operator9:data1]
	signal data_en_0_output_wire                    : std_logic;                     -- data_en_0:output -> [Logical_Bit_Operator10:data1, Logical_Bit_Operator3:data1, cast34:input]
	signal case_statement2_r1_wire                  : std_logic;                     -- Case_Statement2:r1 -> Logical_Bit_Operator3:data0
	signal ctrl_en_0_output_wire                    : std_logic;                     -- ctrl_en_0:output -> [Logical_Bit_Operator4:data0, Logical_Bit_Operator9:data0, cast33:input]
	signal case_statement2_r0_wire                  : std_logic;                     -- Case_Statement2:r0 -> Logical_Bit_Operator4:data1
	signal logical_bit_operator4_result_wire        : std_logic;                     -- Logical_Bit_Operator4:result -> Logical_Bit_Operator5:data0
	signal logical_bit_operator3_result_wire        : std_logic;                     -- Logical_Bit_Operator3:result -> Logical_Bit_Operator5:data1
	signal logical_bit_operator10_result_wire       : std_logic;                     -- Logical_Bit_Operator10:result -> Logical_Bit_Operator6:data1
	signal logical_bit_operator9_result_wire        : std_logic;                     -- Logical_Bit_Operator9:result -> Logical_Bit_Operator6:data0
	signal bus_conversion1_output_wire              : std_logic_vector(1 downto 0);  -- Bus_Conversion1:output -> Multiplexer:sel
	signal delay_output_wire                        : std_logic_vector(23 downto 0); -- Delay:output -> Multiplexer:in0
	signal delay1_output_wire                       : std_logic_vector(23 downto 0); -- Delay1:output -> Multiplexer:in1
	signal delay2_output_wire                       : std_logic_vector(23 downto 0); -- Delay2:output -> Multiplexer:in2
	signal delay3_output_wire                       : std_logic_vector(23 downto 0); -- Delay3:output -> Multiplexer:in3
	signal bus_concatenation_output_wire            : std_logic_vector(1 downto 0);  -- Bus_Concatenation:output -> Multiplexer1:sel
	signal bus_concatenation1_output_wire           : std_logic_vector(1 downto 0);  -- Bus_Concatenation1:output -> Multiplexer2:sel
	signal multiplexer2_result_wire                 : std_logic_vector(24 downto 0); -- Multiplexer2:result -> Multiplexer1:in1
	signal constant18_output_wire                   : std_logic_vector(23 downto 0); -- Constant18:output -> Pipelined_Adder2:datab
	signal pipelined_adder2_result_wire             : std_logic_vector(23 downto 0); -- Pipelined_Adder2:result -> If_Statement7:c
	signal logical_bit_operator5_result_wire        : std_logic;                     -- Logical_Bit_Operator5:result -> sop_0:input
	signal logical_bit_operator6_result_wire        : std_logic;                     -- Logical_Bit_Operator6:result -> eop_0:input
	signal multiplexer1_result_wire                 : std_logic_vector(24 downto 0); -- Multiplexer1:result -> data_0:input
	signal cast29_output_wire                       : std_logic_vector(15 downto 0); -- cast29:output -> Case_Statement1:input
	signal case_statement1_r0_wire                  : std_logic;                     -- Case_Statement1:r0 -> cast30:input
	signal cast30_output_wire                       : std_logic_vector(0 downto 0);  -- cast30:output -> Bus_Concatenation1:a
	signal case_statement1_r1_wire                  : std_logic;                     -- Case_Statement1:r1 -> cast31:input
	signal cast31_output_wire                       : std_logic_vector(0 downto 0);  -- cast31:output -> Bus_Concatenation1:b
	signal cast32_output_wire                       : std_logic_vector(15 downto 0); -- cast32:output -> Case_Statement2:input
	signal cast33_output_wire                       : std_logic_vector(0 downto 0);  -- cast33:output -> Bus_Concatenation:a
	signal cast34_output_wire                       : std_logic_vector(0 downto 0);  -- cast34:output -> Bus_Concatenation:b
	signal constant16_output_wire                   : std_logic_vector(15 downto 0); -- Constant16:output -> cast35:input
	signal cast35_output_wire                       : std_logic_vector(23 downto 0); -- cast35:output -> If_Statement7:b
	signal constant5_output_wire                    : std_logic_vector(23 downto 0); -- Constant5:output -> cast36:input
	signal cast36_output_wire                       : std_logic_vector(24 downto 0); -- cast36:output -> Multiplexer1:in0
	signal multiplexer_result_wire                  : std_logic_vector(23 downto 0); -- Multiplexer:result -> cast37:input
	signal cast37_output_wire                       : std_logic_vector(24 downto 0); -- cast37:output -> Multiplexer1:in2
	signal colorbar_0_output_wire                   : std_logic_vector(23 downto 0); -- colorbar_0:output -> cast38:input
	signal cast38_output_wire                       : std_logic_vector(24 downto 0); -- cast38:output -> Multiplexer2:in0
	signal delay5_output_wire                       : std_logic_vector(23 downto 0); -- Delay5:output -> cast39:input
	signal cast39_output_wire                       : std_logic_vector(24 downto 0); -- cast39:output -> Multiplexer2:in1
	signal pixel_num_0_output_wire                  : std_logic_vector(47 downto 0); -- pixel_num_0:output -> cast40:input
	signal cast40_output_wire                       : std_logic_vector(23 downto 0); -- cast40:output -> Pipelined_Adder2:dataa
	signal clock_0_clock_output_reset               : std_logic;                     -- Clock_0:aclr_out -> [Bus_Concatenation1:aclr, Bus_Concatenation:aclr, Case_Statement1:aclr, Case_Statement2:aclr, Delay1:aclr, Delay2:aclr, Delay3:aclr, Delay5:aclr, Delay:aclr, Multiplexer1:aclr, Multiplexer2:aclr, Multiplexer:aclr, Pipelined_Adder2:aclr]
	signal clock_0_clock_output_clk                 : std_logic;                     -- Clock_0:clock_out -> [Bus_Concatenation1:clock, Bus_Concatenation:clock, Case_Statement1:clock, Case_Statement2:clock, Delay1:clock, Delay2:clock, Delay3:clock, Delay5:clock, Delay:clock, Multiplexer1:clock, Multiplexer2:clock, Multiplexer:clock, Pipelined_Adder2:clock]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	bus_conversion1 : component alt_dspbuilder_cast_GN33BXJAZX
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => counter_0_output_wire,       --  input.wire
			output => bus_conversion1_output_wire  -- output.wire
		);

	pipelined_adder2 : component alt_dspbuilder_pipelined_adder_GNTWZRTG4I
		generic map (
			width    => 24,
			pipeline => 2
		)
		port map (
			clock     => clock_0_clock_output_clk,                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,               --           .reset
			dataa     => cast40_output_wire,                       --      dataa.wire
			datab     => constant18_output_wire,                   --      datab.wire
			result    => pipelined_adder2_result_wire,             --     result.wire
			user_aclr => pipelined_adder2user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder2enavcc_output_wire        --        ena.wire
		);

	pipelined_adder2user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder2user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder2enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder2enavcc_output_wire  -- output.wire
		);

	case_statement1 : component alt_dspbuilder_case_statement_GNWMX2GCN2
		generic map (
			number_outputs => 2,
			hasDefault     => 1,
			pipeline       => 0,
			width          => 16
		)
		port map (
			clock => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset, --           .reset
			input => cast29_output_wire,         --      input.wire
			r0    => case_statement1_r0_wire,    --         r0.wire
			r1    => case_statement1_r1_wire     --         r1.wire
		);

	case_statement2 : component alt_dspbuilder_case_statement_GNFTM45DFU
		generic map (
			number_outputs => 2,
			hasDefault     => 0,
			pipeline       => 0,
			width          => 16
		)
		port map (
			clock => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr  => clock_0_clock_output_reset, --           .reset
			input => cast32_output_wire,         --      input.wire
			r0    => case_statement2_r0_wire,    --         r0.wire
			r1    => case_statement2_r1_wire     --         r1.wire
		);

	multiplexer : component alt_dspbuilder_multiplexer_GNLGLCKYZ5
		generic map (
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0,
			width                  => 24,
			pipeline               => 0,
			number_inputs          => 4
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			sel       => bus_conversion1_output_wire,         --        sel.wire
			result    => multiplexer_result_wire,             --     result.wire
			ena       => multiplexerenavcc_output_wire,       --        ena.wire
			user_aclr => multiplexeruser_aclrgnd_output_wire, --  user_aclr.wire
			in0       => delay_output_wire,                   --        in0.wire
			in1       => delay1_output_wire,                  --        in1.wire
			in2       => delay2_output_wire,                  --        in2.wire
			in3       => delay3_output_wire                   --        in3.wire
		);

	multiplexeruser_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexeruser_aclrgnd_output_wire  -- output.wire
		);

	multiplexerenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexerenavcc_output_wire  -- output.wire
		);

	data_0 : component alt_dspbuilder_port_GNEHYJMBQS
		port map (
			input  => multiplexer1_result_wire, --  input.wire
			output => data                      -- output.wire
		);

	constant7 : component alt_dspbuilder_constant_GNNKZSYI73
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "000000000000000000000000",
			width      => 24
		)
		port map (
			output => constant7_output_wire  -- output.wire
		);

	constant5 : component alt_dspbuilder_constant_GNNKZSYI73
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "000000000000000000000000",
			width      => 24
		)
		port map (
			output => constant5_output_wire  -- output.wire
		);

	bus_concatenation1 : component alt_dspbuilder_bus_concat_GN6E6AAQPZ
		generic map (
			widthB => 1,
			widthA => 1
		)
		port map (
			clock  => clock_0_clock_output_clk,       -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,     --           .reset
			a      => cast30_output_wire,             --          a.wire
			b      => cast31_output_wire,             --          b.wire
			output => bus_concatenation1_output_wire  --     output.wire
		);

	logical_bit_operator6 : component alt_dspbuilder_logical_bit_op_GNUQ2R64DV
		generic map (
			LogicalOp     => "AltOR",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator6_result_wire,  -- result.wire
			data0  => logical_bit_operator9_result_wire,  --  data0.wire
			data1  => logical_bit_operator10_result_wire  --  data1.wire
		);

	logical_bit_operator5 : component alt_dspbuilder_logical_bit_op_GNUQ2R64DV
		generic map (
			LogicalOp     => "AltOR",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator5_result_wire, -- result.wire
			data0  => logical_bit_operator4_result_wire, --  data0.wire
			data1  => logical_bit_operator3_result_wire  --  data1.wire
		);

	ctrl_pak2_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => ctrl_pak2,               --  input.wire
			output => ctrl_pak2_0_output_wire  -- output.wire
		);

	logical_bit_operator4 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator4_result_wire, -- result.wire
			data0  => ctrl_en_0_output_wire,             --  data0.wire
			data1  => case_statement2_r0_wire            --  data1.wire
		);

	ctrl_pak3_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => ctrl_pak3,               --  input.wire
			output => ctrl_pak3_0_output_wire  -- output.wire
		);

	bus_concatenation : component alt_dspbuilder_bus_concat_GN6E6AAQPZ
		generic map (
			widthB => 1,
			widthA => 1
		)
		port map (
			clock  => clock_0_clock_output_clk,      -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset,    --           .reset
			a      => cast33_output_wire,            --          a.wire
			b      => cast34_output_wire,            --          b.wire
			output => bus_concatenation_output_wire  --     output.wire
		);

	ctrl_pak1_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => ctrl_pak1,               --  input.wire
			output => ctrl_pak1_0_output_wire  -- output.wire
		);

	logical_bit_operator9 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator9_result_wire, -- result.wire
			data0  => ctrl_en_0_output_wire,             --  data0.wire
			data1  => if_statement7_true_wire            --  data1.wire
		);

	constant1 : component alt_dspbuilder_constant_GNZEH3JAKA
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "000000000000000000001111",
			width      => 24
		)
		port map (
			output => constant1_output_wire  -- output.wire
		);

	delay : component alt_dspbuilder_delay_GNIYBMGPQQ
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 0,
			BitPattern => "000000000000000000001111",
			width      => 24
		)
		port map (
			input  => constant1_output_wire,      --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay_output_wire,          --     output.wire
			sclr   => delaysclrgnd_output_wire,   --       sclr.wire
			ena    => delayenavcc_output_wire     --        ena.wire
		);

	delaysclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delaysclrgnd_output_wire  -- output.wire
		);

	delayenavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => delayenavcc_output_wire  -- output.wire
		);

	constant16 : component alt_dspbuilder_constant_GNLJWFEWBD
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "0000000000000011",
			width      => 16
		)
		port map (
			output => constant16_output_wire  -- output.wire
		);

	constant18 : component alt_dspbuilder_constant_GNQJ63TWA6
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "000000000000000000000100",
			width      => 24
		)
		port map (
			output => constant18_output_wire  -- output.wire
		);

	logical_bit_operator3 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator3_result_wire, -- result.wire
			data0  => case_statement2_r1_wire,           --  data0.wire
			data1  => data_en_0_output_wire              --  data1.wire
		);

	eop_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => logical_bit_operator6_result_wire, --  input.wire
			output => eop                                -- output.wire
		);

	colorbar_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => colorbar,               --  input.wire
			output => colorbar_0_output_wire  -- output.wire
		);

	if_statement7 : component alt_dspbuilder_if_statement_GNTVBNRAAT
		generic map (
			use_else_output => 0,
			bwr             => 0,
			use_else_input  => 0,
			signed          => 0,
			HDLTYPE         => "STD_LOGIC_VECTOR",
			if_expression   => "(a=b) or (a=c)",
			number_inputs   => 3,
			width           => 24
		)
		port map (
			true => if_statement7_true_wire,      -- true.wire
			a    => counter_0_output_wire,        --    a.wire
			b    => cast35_output_wire,           --    b.wire
			c    => pipelined_adder2_result_wire  --    c.wire
		);

	counter_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => counter,               --  input.wire
			output => counter_0_output_wire  -- output.wire
		);

	delay5 : component alt_dspbuilder_delay_GNNBTO2F3L
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 0,
			BitPattern => "000000000000000000000010",
			width      => 24
		)
		port map (
			input  => constant7_output_wire,      --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay5_output_wire,         --     output.wire
			sclr   => delay5sclrgnd_output_wire,  --       sclr.wire
			ena    => delay5enavcc_output_wire    --        ena.wire
		);

	delay5sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay5sclrgnd_output_wire  -- output.wire
		);

	delay5enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => delay5enavcc_output_wire  -- output.wire
		);

	pixel_num_0 : component alt_dspbuilder_port_GNUJT4YY5I
		port map (
			input  => pixel_num,               --  input.wire
			output => pixel_num_0_output_wire  -- output.wire
		);

	delay3 : component alt_dspbuilder_delay_GNNBTO2F3L
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 0,
			BitPattern => "000000000000000000000010",
			width      => 24
		)
		port map (
			input  => ctrl_pak3_0_output_wire,    --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay3_output_wire,         --     output.wire
			sclr   => delay3sclrgnd_output_wire,  --       sclr.wire
			ena    => delay3enavcc_output_wire    --        ena.wire
		);

	delay3sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay3sclrgnd_output_wire  -- output.wire
		);

	delay3enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => delay3enavcc_output_wire  -- output.wire
		);

	sop_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => logical_bit_operator5_result_wire, --  input.wire
			output => sop                                -- output.wire
		);

	logical_bit_operator10 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator10_result_wire, -- result.wire
			data0  => if_statement7_true_wire,            --  data0.wire
			data1  => data_en_0_output_wire               --  data1.wire
		);

	ctrl_en_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => ctrl_en,               --  input.wire
			output => ctrl_en_0_output_wire  -- output.wire
		);

	multiplexer1 : component alt_dspbuilder_multiplexer_GNHQFFAUXQ
		generic map (
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 0,
			width                  => 25,
			pipeline               => 0,
			number_inputs          => 3
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => bus_concatenation_output_wire,        --        sel.wire
			result    => multiplexer1_result_wire,             --     result.wire
			ena       => multiplexer1enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer1user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => cast36_output_wire,                   --        in0.wire
			in1       => multiplexer2_result_wire,             --        in1.wire
			in2       => cast37_output_wire                    --        in2.wire
		);

	multiplexer1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer1user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer1enavcc_output_wire  -- output.wire
		);

	delay1 : component alt_dspbuilder_delay_GNNBTO2F3L
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 0,
			BitPattern => "000000000000000000000010",
			width      => 24
		)
		port map (
			input  => ctrl_pak1_0_output_wire,    --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay1_output_wire,         --     output.wire
			sclr   => delay1sclrgnd_output_wire,  --       sclr.wire
			ena    => delay1enavcc_output_wire    --        ena.wire
		);

	delay1sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay1sclrgnd_output_wire  -- output.wire
		);

	delay1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => delay1enavcc_output_wire  -- output.wire
		);

	multiplexer2 : component alt_dspbuilder_multiplexer_GN6ODCX3D4
		generic map (
			HDLTYPE                => "STD_LOGIC_VECTOR",
			use_one_hot_select_bus => 1,
			width                  => 25,
			pipeline               => 0,
			number_inputs          => 2
		)
		port map (
			clock     => clock_0_clock_output_clk,             -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,           --           .reset
			sel       => bus_concatenation1_output_wire,       --        sel.wire
			result    => multiplexer2_result_wire,             --     result.wire
			ena       => multiplexer2enavcc_output_wire,       --        ena.wire
			user_aclr => multiplexer2user_aclrgnd_output_wire, --  user_aclr.wire
			in0       => cast38_output_wire,                   --        in0.wire
			in1       => cast39_output_wire                    --        in1.wire
		);

	multiplexer2user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplexer2user_aclrgnd_output_wire  -- output.wire
		);

	multiplexer2enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplexer2enavcc_output_wire  -- output.wire
		);

	delay2 : component alt_dspbuilder_delay_GNVJUPFOX3
		generic map (
			ClockPhase => "1",
			delay      => 1,
			use_init   => 0,
			BitPattern => "000000000000000000000000",
			width      => 24
		)
		port map (
			input  => ctrl_pak2_0_output_wire,    --      input.wire
			clock  => clock_0_clock_output_clk,   -- clock_aclr.clk
			aclr   => clock_0_clock_output_reset, --           .reset
			output => delay2_output_wire,         --     output.wire
			sclr   => delay2sclrgnd_output_wire,  --       sclr.wire
			ena    => delay2enavcc_output_wire    --        ena.wire
		);

	delay2sclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => delay2sclrgnd_output_wire  -- output.wire
		);

	delay2enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => delay2enavcc_output_wire  -- output.wire
		);

	data_en_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => data_en,               --  input.wire
			output => data_en_0_output_wire  -- output.wire
		);

	cast29 : component alt_dspbuilder_cast_GN3ODVPHOL
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => counter_0_output_wire, --  input.wire
			output => cast29_output_wire     -- output.wire
		);

	cast30 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => case_statement1_r0_wire, --  input.wire
			output => cast30_output_wire       -- output.wire
		);

	cast31 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => case_statement1_r1_wire, --  input.wire
			output => cast31_output_wire       -- output.wire
		);

	cast32 : component alt_dspbuilder_cast_GN3ODVPHOL
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => counter_0_output_wire, --  input.wire
			output => cast32_output_wire     -- output.wire
		);

	cast33 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => ctrl_en_0_output_wire, --  input.wire
			output => cast33_output_wire     -- output.wire
		);

	cast34 : component alt_dspbuilder_cast_GN46N4UJ5S
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => data_en_0_output_wire, --  input.wire
			output => cast34_output_wire     -- output.wire
		);

	cast35 : component alt_dspbuilder_cast_GNCPEUNC4M
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant16_output_wire, --  input.wire
			output => cast35_output_wire      -- output.wire
		);

	cast36 : component alt_dspbuilder_cast_GNKDE2NVCC
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => constant5_output_wire, --  input.wire
			output => cast36_output_wire     -- output.wire
		);

	cast37 : component alt_dspbuilder_cast_GNKDE2NVCC
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplexer_result_wire, --  input.wire
			output => cast37_output_wire       -- output.wire
		);

	cast38 : component alt_dspbuilder_cast_GNCCZ56SYK
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => colorbar_0_output_wire, --  input.wire
			output => cast38_output_wire      -- output.wire
		);

	cast39 : component alt_dspbuilder_cast_GNKDE2NVCC
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => delay5_output_wire, --  input.wire
			output => cast39_output_wire  -- output.wire
		);

	cast40 : component alt_dspbuilder_cast_GNKIWLRTQI
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => pixel_num_0_output_wire, --  input.wire
			output => cast40_output_wire       -- output.wire
		);

end architecture rtl; -- of Test_Pattern_Generator_GN_Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT
