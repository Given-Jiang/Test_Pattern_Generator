-- Test_Pattern_Generator_GN_Test_Pattern_Generator_MAIN_CTRL.vhd

-- Generated using ACDS version 13.1 162 at 2015.02.27.10:05:29

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Test_Pattern_Generator_GN_Test_Pattern_Generator_MAIN_CTRL is
	port (
		eop       : out std_logic;                                        --       eop.wire
		counter_1 : out std_logic_vector(23 downto 0);                    -- counter_1.wire
		colorbar  : in  std_logic_vector(23 downto 0) := (others => '0'); --  colorbar.wire
		data      : out std_logic_vector(24 downto 0);                    --      data.wire
		col       : in  std_logic_vector(31 downto 0) := (others => '0'); --       col.wire
		ctrl_pak3 : in  std_logic_vector(23 downto 0) := (others => '0'); -- ctrl_pak3.wire
		ctrl_pak2 : in  std_logic_vector(23 downto 0) := (others => '0'); -- ctrl_pak2.wire
		data_en   : out std_logic;                                        --   data_en.wire
		ctrl_en   : out std_logic;                                        --   ctrl_en.wire
		Clock     : in  std_logic                     := '0';             --     Clock.clk
		aclr      : in  std_logic                     := '0';             --          .reset
		row       : in  std_logic_vector(31 downto 0) := (others => '0'); --       row.wire
		ctrl_pak1 : in  std_logic_vector(23 downto 0) := (others => '0'); -- ctrl_pak1.wire
		check_en  : out std_logic;                                        --  check_en.wire
		sop       : out std_logic;                                        --       sop.wire
		ready     : in  std_logic                     := '0'              --     ready.wire
	);
end entity Test_Pattern_Generator_GN_Test_Pattern_Generator_MAIN_CTRL;

architecture rtl of Test_Pattern_Generator_GN_Test_Pattern_Generator_MAIN_CTRL is
	component alt_dspbuilder_clock_GNQFU4PUDH is
		port (
			aclr      : in  std_logic := 'X'; -- reset
			aclr_n    : in  std_logic := 'X'; -- reset_n
			aclr_out  : out std_logic;        -- reset
			clock     : in  std_logic := 'X'; -- clk
			clock_out : out std_logic         -- clk
		);
	end component alt_dspbuilder_clock_GNQFU4PUDH;

	component alt_dspbuilder_port_GNEPKLLZKY is
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(31 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNEPKLLZKY;

	component alt_dspbuilder_port_GNOC3SGKQJ is
		port (
			input  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNOC3SGKQJ;

	component alt_dspbuilder_pipelined_adder_GNTWZRTG4I is
		generic (
			width    : natural := 0;
			pipeline : integer := 0
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			add_sub   : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cout      : out std_logic;                                             -- wire
			dataa     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			datab     : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			result    : out std_logic_vector(width-1 downto 0);                    -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_pipelined_adder_GNTWZRTG4I;

	component alt_dspbuilder_gnd_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_gnd_GN;

	component alt_dspbuilder_vcc_GN is
		port (
			output : out std_logic   -- wire
		);
	end component alt_dspbuilder_vcc_GN;

	component alt_dspbuilder_port_GNEHYJMBQS is
		port (
			input  : in  std_logic_vector(24 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(24 downto 0)                     -- wire
		);
	end component alt_dspbuilder_port_GNEHYJMBQS;

	component alt_dspbuilder_if_statement_GNIV4UP6ZO is
		generic (
			use_else_output : natural := 0;
			bwr             : natural := 0;
			use_else_input  : natural := 0;
			signed          : natural := 1;
			HDLTYPE         : string  := "STD_LOGIC_VECTOR";
			if_expression   : string  := "a";
			number_inputs   : integer := 1;
			width           : natural := 8
		);
		port (
			true : out std_logic;                                        -- wire
			a    : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			b    : in  std_logic_vector(23 downto 0) := (others => 'X')  -- wire
		);
	end component alt_dspbuilder_if_statement_GNIV4UP6ZO;

	component alt_dspbuilder_counter_GNKAA2ZBZG is
		generic (
			use_usr_aclr : string  := "false";
			use_ena      : string  := "false";
			use_cin      : string  := "false";
			use_sset     : string  := "false";
			ndirection   : natural := 1;
			svalue       : string  := "0";
			use_sload    : string  := "false";
			use_sclr     : string  := "false";
			use_cout     : string  := "false";
			modulus      : integer := 256;
			use_cnt_ena  : string  := "false";
			width        : natural := 8;
			use_aset     : string  := "false";
			use_aload    : string  := "false";
			avalue       : string  := "0"
		);
		port (
			aclr      : in  std_logic                          := 'X';             -- clk
			aload     : in  std_logic                          := 'X';             -- wire
			aset      : in  std_logic                          := 'X';             -- wire
			cin       : in  std_logic                          := 'X';             -- wire
			clock     : in  std_logic                          := 'X';             -- clk
			cnt_ena   : in  std_logic                          := 'X';             -- wire
			cout      : out std_logic;                                             -- wire
			data      : in  std_logic_vector(width-1 downto 0) := (others => 'X'); -- wire
			direction : in  std_logic                          := 'X';             -- wire
			ena       : in  std_logic                          := 'X';             -- wire
			q         : out std_logic_vector(width-1 downto 0);                    -- wire
			sclr      : in  std_logic                          := 'X';             -- wire
			sload     : in  std_logic                          := 'X';             -- wire
			sset      : in  std_logic                          := 'X';             -- wire
			user_aclr : in  std_logic                          := 'X'              -- wire
		);
	end component alt_dspbuilder_counter_GNKAA2ZBZG;

	component alt_dspbuilder_constant_GNQJ63TWA6 is
		generic (
			HDLTYPE    : string  := "STD_LOGIC_VECTOR";
			BitPattern : string  := "0000";
			width      : natural := 4
		);
		port (
			output : out std_logic_vector(23 downto 0)   -- wire
		);
	end component alt_dspbuilder_constant_GNQJ63TWA6;

	component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'; -- wire
			data1  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V;

	component alt_dspbuilder_port_GN37ALZBS4 is
		port (
			input  : in  std_logic := 'X'; -- wire
			output : out std_logic         -- wire
		);
	end component alt_dspbuilder_port_GN37ALZBS4;

	component Test_Pattern_Generator_GN_Test_Pattern_Generator_MAIN_CTRL_CTRL_TOP is
		port (
			Clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X';             -- reset
			check_en  : out std_logic;                                        -- wire
			pixel_num : in  std_logic_vector(47 downto 0) := (others => 'X'); -- wire
			ready     : in  std_logic                     := 'X';             -- wire
			data_en   : out std_logic;                                        -- wire
			counter   : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			ctrl_en   : out std_logic                                         -- wire
		);
	end component Test_Pattern_Generator_GN_Test_Pattern_Generator_MAIN_CTRL_CTRL_TOP;

	component alt_dspbuilder_multiplier_GNEIWYOKUR is
		generic (
			DEDICATED_MULTIPLIER_CIRCUITRY : string  := "AUTO";
			Signed                         : natural := 0;
			OutputMsb                      : integer := 8;
			aWidth                         : natural := 8;
			bWidth                         : natural := 8;
			OutputLsb                      : integer := 0;
			pipeline                       : integer := 0
		);
		port (
			aclr      : in  std_logic                                          := 'X';             -- clk
			clock     : in  std_logic                                          := 'X';             -- clk
			dataa     : in  std_logic_vector(aWidth-1 downto 0)                := (others => 'X'); -- wire
			datab     : in  std_logic_vector(bWidth-1 downto 0)                := (others => 'X'); -- wire
			ena       : in  std_logic                                          := 'X';             -- wire
			result    : out std_logic_vector(OutputMsb-OutputLsb+1-1 downto 0);                    -- wire
			user_aclr : in  std_logic                                          := 'X'              -- wire
		);
	end component alt_dspbuilder_multiplier_GNEIWYOKUR;

	component Test_Pattern_Generator_GN_Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT is
		port (
			sop       : out std_logic;                                        -- wire
			pixel_num : in  std_logic_vector(47 downto 0) := (others => 'X'); -- wire
			ctrl_en   : in  std_logic                     := 'X';             -- wire
			counter   : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			ctrl_pak1 : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			colorbar  : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			data      : out std_logic_vector(24 downto 0);                    -- wire
			data_en   : in  std_logic                     := 'X';             -- wire
			ctrl_pak2 : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			eop       : out std_logic;                                        -- wire
			ctrl_pak3 : in  std_logic_vector(23 downto 0) := (others => 'X'); -- wire
			Clock     : in  std_logic                     := 'X';             -- clk
			aclr      : in  std_logic                     := 'X'              -- reset
		);
	end component Test_Pattern_Generator_GN_Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT;

	component alt_dspbuilder_logical_bit_op_GNUQ2R64DV is
		generic (
			LogicalOp     : string   := "AltAND";
			number_inputs : positive := 2
		);
		port (
			result : out std_logic;        -- wire
			data0  : in  std_logic := 'X'; -- wire
			data1  : in  std_logic := 'X'  -- wire
		);
	end component alt_dspbuilder_logical_bit_op_GNUQ2R64DV;

	component alt_dspbuilder_cast_GN7PRGDOVA is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GN7PRGDOVA;

	component alt_dspbuilder_cast_GNKIWLRTQI is
		generic (
			round    : natural := 0;
			saturate : natural := 0
		);
		port (
			input  : in  std_logic_vector(47 downto 0) := (others => 'X'); -- wire
			output : out std_logic_vector(23 downto 0)                     -- wire
		);
	end component alt_dspbuilder_cast_GNKIWLRTQI;

	signal pipelined_adder5user_aclrgnd_output_wire                  : std_logic;                     -- Pipelined_Adder5user_aclrGND:output -> Pipelined_Adder5:user_aclr
	signal pipelined_adder5enavcc_output_wire                        : std_logic;                     -- Pipelined_Adder5enaVCC:output -> Pipelined_Adder5:ena
	signal multiplier1user_aclrgnd_output_wire                       : std_logic;                     -- Multiplier1user_aclrGND:output -> Multiplier1:user_aclr
	signal multiplier1enavcc_output_wire                             : std_logic;                     -- Multiplier1enaVCC:output -> Multiplier1:ena
	signal ready_0_output_wire                                       : std_logic;                     -- ready_0:output -> Test_Pattern_Generator_MAIN_CTRL_CTRL_TOP_0:ready
	signal counter_q_wire                                            : std_logic_vector(23 downto 0); -- Counter:q -> [If_Statement4:a, Test_Pattern_Generator_MAIN_CTRL_CTRL_TOP_0:counter, Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT_0:counter, counter_1_0:input]
	signal test_pattern_generator_main_ctrl_ctrl_top_0_ctrl_en_wire  : std_logic;                     -- Test_Pattern_Generator_MAIN_CTRL_CTRL_TOP_0:ctrl_en -> [Logical_Bit_Operator1:data0, Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT_0:ctrl_en, ctrl_en_0:input]
	signal test_pattern_generator_main_ctrl_ctrl_top_0_data_en_wire  : std_logic;                     -- Test_Pattern_Generator_MAIN_CTRL_CTRL_TOP_0:data_en -> [Logical_Bit_Operator11:data0, Logical_Bit_Operator1:data1, Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT_0:data_en, data_en_0:input]
	signal logical_bit_operator1_result_wire                         : std_logic;                     -- Logical_Bit_Operator1:result -> Counter:cnt_ena
	signal if_statement4_true_wire                                   : std_logic;                     -- If_Statement4:true -> Logical_Bit_Operator11:data1
	signal logical_bit_operator11_result_wire                        : std_logic;                     -- Logical_Bit_Operator11:result -> Counter:sclr
	signal multiplier1_result_wire                                   : std_logic_vector(47 downto 0); -- Multiplier1:result -> [Test_Pattern_Generator_MAIN_CTRL_CTRL_TOP_0:pixel_num, Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT_0:pixel_num, cast43:input]
	signal constant4_output_wire                                     : std_logic_vector(23 downto 0); -- Constant4:output -> Pipelined_Adder5:datab
	signal pipelined_adder5_result_wire                              : std_logic_vector(23 downto 0); -- Pipelined_Adder5:result -> If_Statement4:b
	signal ctrl_pak1_0_output_wire                                   : std_logic_vector(23 downto 0); -- ctrl_pak1_0:output -> Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT_0:ctrl_pak1
	signal ctrl_pak2_0_output_wire                                   : std_logic_vector(23 downto 0); -- ctrl_pak2_0:output -> Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT_0:ctrl_pak2
	signal ctrl_pak3_0_output_wire                                   : std_logic_vector(23 downto 0); -- ctrl_pak3_0:output -> Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT_0:ctrl_pak3
	signal colorbar_0_output_wire                                    : std_logic_vector(23 downto 0); -- colorbar_0:output -> Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT_0:colorbar
	signal test_pattern_generator_main_ctrl_signal_out_0_data_wire   : std_logic_vector(24 downto 0); -- Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT_0:data -> data_0:input
	signal test_pattern_generator_main_ctrl_signal_out_0_sop_wire    : std_logic;                     -- Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT_0:sop -> sop_0:input
	signal test_pattern_generator_main_ctrl_signal_out_0_eop_wire    : std_logic;                     -- Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT_0:eop -> eop_0:input
	signal test_pattern_generator_main_ctrl_ctrl_top_0_check_en_wire : std_logic;                     -- Test_Pattern_Generator_MAIN_CTRL_CTRL_TOP_0:check_en -> check_en_0:input
	signal col_0_output_wire                                         : std_logic_vector(31 downto 0); -- col_0:output -> cast41:input
	signal cast41_output_wire                                        : std_logic_vector(23 downto 0); -- cast41:output -> Multiplier1:dataa
	signal row_0_output_wire                                         : std_logic_vector(31 downto 0); -- row_0:output -> cast42:input
	signal cast42_output_wire                                        : std_logic_vector(23 downto 0); -- cast42:output -> Multiplier1:datab
	signal cast43_output_wire                                        : std_logic_vector(23 downto 0); -- cast43:output -> Pipelined_Adder5:dataa
	signal clock_0_clock_output_reset                                : std_logic;                     -- Clock_0:aclr_out -> [Counter:aclr, Multiplier1:aclr, Pipelined_Adder5:aclr, Test_Pattern_Generator_MAIN_CTRL_CTRL_TOP_0:aclr, Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT_0:aclr]
	signal clock_0_clock_output_clk                                  : std_logic;                     -- Clock_0:clock_out -> [Counter:clock, Multiplier1:clock, Pipelined_Adder5:clock, Test_Pattern_Generator_MAIN_CTRL_CTRL_TOP_0:Clock, Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT_0:Clock]

begin

	clock_0 : component alt_dspbuilder_clock_GNQFU4PUDH
		port map (
			clock_out => clock_0_clock_output_clk,   -- clock_output.clk
			aclr_out  => clock_0_clock_output_reset, --             .reset
			clock     => Clock,                      --        clock.clk
			aclr      => aclr                        --             .reset
		);

	col_0 : component alt_dspbuilder_port_GNEPKLLZKY
		port map (
			input  => col,               --  input.wire
			output => col_0_output_wire  -- output.wire
		);

	counter_1_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => counter_q_wire, --  input.wire
			output => counter_1       -- output.wire
		);

	colorbar_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => colorbar,               --  input.wire
			output => colorbar_0_output_wire  -- output.wire
		);

	pipelined_adder5 : component alt_dspbuilder_pipelined_adder_GNTWZRTG4I
		generic map (
			width    => 24,
			pipeline => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,                 -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,               --           .reset
			dataa     => cast43_output_wire,                       --      dataa.wire
			datab     => constant4_output_wire,                    --      datab.wire
			result    => pipelined_adder5_result_wire,             --     result.wire
			user_aclr => pipelined_adder5user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => pipelined_adder5enavcc_output_wire        --        ena.wire
		);

	pipelined_adder5user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => pipelined_adder5user_aclrgnd_output_wire  -- output.wire
		);

	pipelined_adder5enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => pipelined_adder5enavcc_output_wire  -- output.wire
		);

	data_0 : component alt_dspbuilder_port_GNEHYJMBQS
		port map (
			input  => test_pattern_generator_main_ctrl_signal_out_0_data_wire, --  input.wire
			output => data                                                     -- output.wire
		);

	if_statement4 : component alt_dspbuilder_if_statement_GNIV4UP6ZO
		generic map (
			use_else_output => 0,
			bwr             => 0,
			use_else_input  => 0,
			signed          => 0,
			HDLTYPE         => "STD_LOGIC_VECTOR",
			if_expression   => "a=b",
			number_inputs   => 2,
			width           => 24
		)
		port map (
			true => if_statement4_true_wire,      -- true.wire
			a    => counter_q_wire,               --    a.wire
			b    => pipelined_adder5_result_wire  --    b.wire
		);

	counter : component alt_dspbuilder_counter_GNKAA2ZBZG
		generic map (
			use_usr_aclr => "false",
			use_ena      => "false",
			use_cin      => "false",
			use_sset     => "false",
			ndirection   => 1,
			svalue       => "1",
			use_sload    => "false",
			use_sclr     => "true",
			use_cout     => "false",
			modulus      => 8388608,
			use_cnt_ena  => "true",
			width        => 24,
			use_aset     => "false",
			use_aload    => "false",
			avalue       => "0"
		)
		port map (
			clock   => clock_0_clock_output_clk,           -- clock_aclr.clk
			aclr    => clock_0_clock_output_reset,         --           .reset
			cnt_ena => logical_bit_operator1_result_wire,  --    cnt_ena.wire
			sclr    => logical_bit_operator11_result_wire, --       sclr.wire
			q       => counter_q_wire,                     --          q.wire
			cout    => open                                --       cout.wire
		);

	constant4 : component alt_dspbuilder_constant_GNQJ63TWA6
		generic map (
			HDLTYPE    => "STD_LOGIC_VECTOR",
			BitPattern => "000000000000000000000100",
			width      => 24
		)
		port map (
			output => constant4_output_wire  -- output.wire
		);

	logical_bit_operator11 : component alt_dspbuilder_logical_bit_op_GNA5ZFEL7V
		generic map (
			LogicalOp     => "AltAND",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator11_result_wire,                       -- result.wire
			data0  => test_pattern_generator_main_ctrl_ctrl_top_0_data_en_wire, --  data0.wire
			data1  => if_statement4_true_wire                                   --  data1.wire
		);

	sop_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => test_pattern_generator_main_ctrl_signal_out_0_sop_wire, --  input.wire
			output => sop                                                     -- output.wire
		);

	ready_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => ready,               --  input.wire
			output => ready_0_output_wire  -- output.wire
		);

	row_0 : component alt_dspbuilder_port_GNEPKLLZKY
		port map (
			input  => row,               --  input.wire
			output => row_0_output_wire  -- output.wire
		);

	test_pattern_generator_main_ctrl_ctrl_top_0 : component Test_Pattern_Generator_GN_Test_Pattern_Generator_MAIN_CTRL_CTRL_TOP
		port map (
			Clock     => clock_0_clock_output_clk,                                  --     Clock.clk
			aclr      => clock_0_clock_output_reset,                                --          .reset
			check_en  => test_pattern_generator_main_ctrl_ctrl_top_0_check_en_wire, --  check_en.wire
			pixel_num => multiplier1_result_wire,                                   -- pixel_num.wire
			ready     => ready_0_output_wire,                                       --     ready.wire
			data_en   => test_pattern_generator_main_ctrl_ctrl_top_0_data_en_wire,  --   data_en.wire
			counter   => counter_q_wire,                                            --   counter.wire
			ctrl_en   => test_pattern_generator_main_ctrl_ctrl_top_0_ctrl_en_wire   --   ctrl_en.wire
		);

	ctrl_en_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => test_pattern_generator_main_ctrl_ctrl_top_0_ctrl_en_wire, --  input.wire
			output => ctrl_en                                                   -- output.wire
		);

	ctrl_pak2_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => ctrl_pak2,               --  input.wire
			output => ctrl_pak2_0_output_wire  -- output.wire
		);

	ctrl_pak3_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => ctrl_pak3,               --  input.wire
			output => ctrl_pak3_0_output_wire  -- output.wire
		);

	ctrl_pak1_0 : component alt_dspbuilder_port_GNOC3SGKQJ
		port map (
			input  => ctrl_pak1,               --  input.wire
			output => ctrl_pak1_0_output_wire  -- output.wire
		);

	data_en_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => test_pattern_generator_main_ctrl_ctrl_top_0_data_en_wire, --  input.wire
			output => data_en                                                   -- output.wire
		);

	multiplier1 : component alt_dspbuilder_multiplier_GNEIWYOKUR
		generic map (
			DEDICATED_MULTIPLIER_CIRCUITRY => "YES",
			Signed                         => 0,
			OutputMsb                      => 47,
			aWidth                         => 24,
			bWidth                         => 24,
			OutputLsb                      => 0,
			pipeline                       => 0
		)
		port map (
			clock     => clock_0_clock_output_clk,            -- clock_aclr.clk
			aclr      => clock_0_clock_output_reset,          --           .reset
			dataa     => cast41_output_wire,                  --      dataa.wire
			datab     => cast42_output_wire,                  --      datab.wire
			result    => multiplier1_result_wire,             --     result.wire
			user_aclr => multiplier1user_aclrgnd_output_wire, --  user_aclr.wire
			ena       => multiplier1enavcc_output_wire        --        ena.wire
		);

	multiplier1user_aclrgnd : component alt_dspbuilder_gnd_GN
		port map (
			output => multiplier1user_aclrgnd_output_wire  -- output.wire
		);

	multiplier1enavcc : component alt_dspbuilder_vcc_GN
		port map (
			output => multiplier1enavcc_output_wire  -- output.wire
		);

	test_pattern_generator_main_ctrl_signal_out_0 : component Test_Pattern_Generator_GN_Test_Pattern_Generator_MAIN_CTRL_SIGNAL_OUT
		port map (
			sop       => test_pattern_generator_main_ctrl_signal_out_0_sop_wire,   --       sop.wire
			pixel_num => multiplier1_result_wire,                                  -- pixel_num.wire
			ctrl_en   => test_pattern_generator_main_ctrl_ctrl_top_0_ctrl_en_wire, --   ctrl_en.wire
			counter   => counter_q_wire,                                           --   counter.wire
			ctrl_pak1 => ctrl_pak1_0_output_wire,                                  -- ctrl_pak1.wire
			colorbar  => colorbar_0_output_wire,                                   --  colorbar.wire
			data      => test_pattern_generator_main_ctrl_signal_out_0_data_wire,  --      data.wire
			data_en   => test_pattern_generator_main_ctrl_ctrl_top_0_data_en_wire, --   data_en.wire
			ctrl_pak2 => ctrl_pak2_0_output_wire,                                  -- ctrl_pak2.wire
			eop       => test_pattern_generator_main_ctrl_signal_out_0_eop_wire,   --       eop.wire
			ctrl_pak3 => ctrl_pak3_0_output_wire,                                  -- ctrl_pak3.wire
			Clock     => clock_0_clock_output_clk,                                 --     Clock.clk
			aclr      => clock_0_clock_output_reset                                --          .reset
		);

	check_en_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => test_pattern_generator_main_ctrl_ctrl_top_0_check_en_wire, --  input.wire
			output => check_en                                                   -- output.wire
		);

	eop_0 : component alt_dspbuilder_port_GN37ALZBS4
		port map (
			input  => test_pattern_generator_main_ctrl_signal_out_0_eop_wire, --  input.wire
			output => eop                                                     -- output.wire
		);

	logical_bit_operator1 : component alt_dspbuilder_logical_bit_op_GNUQ2R64DV
		generic map (
			LogicalOp     => "AltOR",
			number_inputs => 2
		)
		port map (
			result => logical_bit_operator1_result_wire,                        -- result.wire
			data0  => test_pattern_generator_main_ctrl_ctrl_top_0_ctrl_en_wire, --  data0.wire
			data1  => test_pattern_generator_main_ctrl_ctrl_top_0_data_en_wire  --  data1.wire
		);

	cast41 : component alt_dspbuilder_cast_GN7PRGDOVA
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => col_0_output_wire,  --  input.wire
			output => cast41_output_wire  -- output.wire
		);

	cast42 : component alt_dspbuilder_cast_GN7PRGDOVA
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => row_0_output_wire,  --  input.wire
			output => cast42_output_wire  -- output.wire
		);

	cast43 : component alt_dspbuilder_cast_GNKIWLRTQI
		generic map (
			round    => 0,
			saturate => 0
		)
		port map (
			input  => multiplier1_result_wire, --  input.wire
			output => cast43_output_wire       -- output.wire
		);

end architecture rtl; -- of Test_Pattern_Generator_GN_Test_Pattern_Generator_MAIN_CTRL
